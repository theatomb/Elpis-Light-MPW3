VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO custom_sram
  CLASS BLOCK ;
  FOREIGN custom_sram ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1500.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 1496.000 23.370 1500.000 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 1496.000 392.290 1500.000 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 670.520 1200.000 671.120 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.200 4.000 637.800 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 0.000 756.610 4.000 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 749.400 1200.000 750.000 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.080 4.000 937.680 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 1496.000 669.210 1500.000 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 1496.000 761.670 1500.000 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 828.960 1200.000 829.560 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 1496.000 115.370 1500.000 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 1496.000 161.830 1500.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 197.240 1200.000 197.840 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 355.000 1200.000 355.600 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 1496.000 300.290 1500.000 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 512.760 1200.000 513.360 ;
    END
  END a[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END clk
  PIN csb0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END csb0_to_sram
  PIN d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END d[0]
  PIN d[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END d[10]
  PIN d[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END d[11]
  PIN d[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 1496.000 438.750 1500.000 ;
    END
  END d[12]
  PIN d[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END d[13]
  PIN d[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END d[14]
  PIN d[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 1496.000 530.750 1500.000 ;
    END
  END d[15]
  PIN d[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.730 0.000 913.010 4.000 ;
    END
  END d[16]
  PIN d[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END d[17]
  PIN d[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 0.000 964.990 4.000 ;
    END
  END d[18]
  PIN d[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 0.000 1017.430 4.000 ;
    END
  END d[19]
  PIN d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END d[1]
  PIN d[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 1496.000 854.130 1500.000 ;
    END
  END d[20]
  PIN d[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 907.840 1200.000 908.440 ;
    END
  END d[21]
  PIN d[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 986.720 1200.000 987.320 ;
    END
  END d[22]
  PIN d[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.160 4.000 1162.760 ;
    END
  END d[23]
  PIN d[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1144.480 1200.000 1145.080 ;
    END
  END d[24]
  PIN d[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 1496.000 1038.590 1500.000 ;
    END
  END d[25]
  PIN d[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1302.240 1200.000 1302.840 ;
    END
  END d[26]
  PIN d[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1312.440 4.000 1313.040 ;
    END
  END d[27]
  PIN d[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END d[28]
  PIN d[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1381.120 1200.000 1381.720 ;
    END
  END d[29]
  PIN d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END d[2]
  PIN d[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.570 0.000 1121.850 4.000 ;
    END
  END d[30]
  PIN d[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.550 0.000 1173.830 4.000 ;
    END
  END d[31]
  PIN d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END d[3]
  PIN d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END d[4]
  PIN d[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END d[5]
  PIN d[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 276.120 1200.000 276.720 ;
    END
  END d[6]
  PIN d[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 1496.000 253.830 1500.000 ;
    END
  END d[7]
  PIN d[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 433.880 1200.000 434.480 ;
    END
  END d[8]
  PIN d[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 1496.000 346.290 1500.000 ;
    END
  END d[9]
  PIN q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 1496.000 69.370 1500.000 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END q[11]
  PIN q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 1496.000 484.750 1500.000 ;
    END
  END q[12]
  PIN q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END q[13]
  PIN q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END q[14]
  PIN q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 1496.000 577.210 1500.000 ;
    END
  END q[15]
  PIN q[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 1496.000 623.210 1500.000 ;
    END
  END q[16]
  PIN q[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 1496.000 715.670 1500.000 ;
    END
  END q[17]
  PIN q[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 1496.000 807.670 1500.000 ;
    END
  END q[18]
  PIN q[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1087.360 4.000 1087.960 ;
    END
  END q[19]
  PIN q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 39.480 1200.000 40.080 ;
    END
  END q[1]
  PIN q[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1496.000 900.130 1500.000 ;
    END
  END q[20]
  PIN q[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.850 1496.000 946.130 1500.000 ;
    END
  END q[21]
  PIN q[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1065.600 1200.000 1066.200 ;
    END
  END q[22]
  PIN q[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 1496.000 992.590 1500.000 ;
    END
  END q[23]
  PIN q[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.960 4.000 1237.560 ;
    END
  END q[24]
  PIN q[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1223.360 1200.000 1223.960 ;
    END
  END q[25]
  PIN q[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 1496.000 1084.590 1500.000 ;
    END
  END q[26]
  PIN q[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1387.240 4.000 1387.840 ;
    END
  END q[27]
  PIN q[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.130 0.000 1069.410 4.000 ;
    END
  END q[28]
  PIN q[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1460.000 1200.000 1460.600 ;
    END
  END q[29]
  PIN q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END q[2]
  PIN q[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.770 1496.000 1131.050 1500.000 ;
    END
  END q[30]
  PIN q[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 1496.000 1177.050 1500.000 ;
    END
  END q[31]
  PIN q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 118.360 1200.000 118.960 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 1496.000 207.830 1500.000 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 591.640 1200.000 592.240 ;
    END
  END q[9]
  PIN spare_wen0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
  END vssd1
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END we
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1195.395 1487.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 1195.455 1488.080 ;
      LAYER met2 ;
        RECT 6.990 1495.720 22.810 1496.000 ;
        RECT 23.650 1495.720 68.810 1496.000 ;
        RECT 69.650 1495.720 114.810 1496.000 ;
        RECT 115.650 1495.720 161.270 1496.000 ;
        RECT 162.110 1495.720 207.270 1496.000 ;
        RECT 208.110 1495.720 253.270 1496.000 ;
        RECT 254.110 1495.720 299.730 1496.000 ;
        RECT 300.570 1495.720 345.730 1496.000 ;
        RECT 346.570 1495.720 391.730 1496.000 ;
        RECT 392.570 1495.720 438.190 1496.000 ;
        RECT 439.030 1495.720 484.190 1496.000 ;
        RECT 485.030 1495.720 530.190 1496.000 ;
        RECT 531.030 1495.720 576.650 1496.000 ;
        RECT 577.490 1495.720 622.650 1496.000 ;
        RECT 623.490 1495.720 668.650 1496.000 ;
        RECT 669.490 1495.720 715.110 1496.000 ;
        RECT 715.950 1495.720 761.110 1496.000 ;
        RECT 761.950 1495.720 807.110 1496.000 ;
        RECT 807.950 1495.720 853.570 1496.000 ;
        RECT 854.410 1495.720 899.570 1496.000 ;
        RECT 900.410 1495.720 945.570 1496.000 ;
        RECT 946.410 1495.720 992.030 1496.000 ;
        RECT 992.870 1495.720 1038.030 1496.000 ;
        RECT 1038.870 1495.720 1084.030 1496.000 ;
        RECT 1084.870 1495.720 1130.490 1496.000 ;
        RECT 1131.330 1495.720 1176.490 1496.000 ;
        RECT 1177.330 1495.720 1190.850 1496.000 ;
        RECT 6.990 4.280 1190.850 1495.720 ;
        RECT 6.990 3.670 25.570 4.280 ;
        RECT 26.410 3.670 77.550 4.280 ;
        RECT 78.390 3.670 129.530 4.280 ;
        RECT 130.370 3.670 181.970 4.280 ;
        RECT 182.810 3.670 233.950 4.280 ;
        RECT 234.790 3.670 286.390 4.280 ;
        RECT 287.230 3.670 338.370 4.280 ;
        RECT 339.210 3.670 390.810 4.280 ;
        RECT 391.650 3.670 442.790 4.280 ;
        RECT 443.630 3.670 494.770 4.280 ;
        RECT 495.610 3.670 547.210 4.280 ;
        RECT 548.050 3.670 599.190 4.280 ;
        RECT 600.030 3.670 651.630 4.280 ;
        RECT 652.470 3.670 703.610 4.280 ;
        RECT 704.450 3.670 756.050 4.280 ;
        RECT 756.890 3.670 808.030 4.280 ;
        RECT 808.870 3.670 860.010 4.280 ;
        RECT 860.850 3.670 912.450 4.280 ;
        RECT 913.290 3.670 964.430 4.280 ;
        RECT 965.270 3.670 1016.870 4.280 ;
        RECT 1017.710 3.670 1068.850 4.280 ;
        RECT 1069.690 3.670 1121.290 4.280 ;
        RECT 1122.130 3.670 1173.270 4.280 ;
        RECT 1174.110 3.670 1190.850 4.280 ;
      LAYER met3 ;
        RECT 4.000 1463.040 1196.000 1488.005 ;
        RECT 4.400 1461.640 1196.000 1463.040 ;
        RECT 4.000 1461.000 1196.000 1461.640 ;
        RECT 4.000 1459.600 1195.600 1461.000 ;
        RECT 4.000 1388.240 1196.000 1459.600 ;
        RECT 4.400 1386.840 1196.000 1388.240 ;
        RECT 4.000 1382.120 1196.000 1386.840 ;
        RECT 4.000 1380.720 1195.600 1382.120 ;
        RECT 4.000 1313.440 1196.000 1380.720 ;
        RECT 4.400 1312.040 1196.000 1313.440 ;
        RECT 4.000 1303.240 1196.000 1312.040 ;
        RECT 4.000 1301.840 1195.600 1303.240 ;
        RECT 4.000 1237.960 1196.000 1301.840 ;
        RECT 4.400 1236.560 1196.000 1237.960 ;
        RECT 4.000 1224.360 1196.000 1236.560 ;
        RECT 4.000 1222.960 1195.600 1224.360 ;
        RECT 4.000 1163.160 1196.000 1222.960 ;
        RECT 4.400 1161.760 1196.000 1163.160 ;
        RECT 4.000 1145.480 1196.000 1161.760 ;
        RECT 4.000 1144.080 1195.600 1145.480 ;
        RECT 4.000 1088.360 1196.000 1144.080 ;
        RECT 4.400 1086.960 1196.000 1088.360 ;
        RECT 4.000 1066.600 1196.000 1086.960 ;
        RECT 4.000 1065.200 1195.600 1066.600 ;
        RECT 4.000 1012.880 1196.000 1065.200 ;
        RECT 4.400 1011.480 1196.000 1012.880 ;
        RECT 4.000 987.720 1196.000 1011.480 ;
        RECT 4.000 986.320 1195.600 987.720 ;
        RECT 4.000 938.080 1196.000 986.320 ;
        RECT 4.400 936.680 1196.000 938.080 ;
        RECT 4.000 908.840 1196.000 936.680 ;
        RECT 4.000 907.440 1195.600 908.840 ;
        RECT 4.000 863.280 1196.000 907.440 ;
        RECT 4.400 861.880 1196.000 863.280 ;
        RECT 4.000 829.960 1196.000 861.880 ;
        RECT 4.000 828.560 1195.600 829.960 ;
        RECT 4.000 788.480 1196.000 828.560 ;
        RECT 4.400 787.080 1196.000 788.480 ;
        RECT 4.000 750.400 1196.000 787.080 ;
        RECT 4.000 749.000 1195.600 750.400 ;
        RECT 4.000 713.000 1196.000 749.000 ;
        RECT 4.400 711.600 1196.000 713.000 ;
        RECT 4.000 671.520 1196.000 711.600 ;
        RECT 4.000 670.120 1195.600 671.520 ;
        RECT 4.000 638.200 1196.000 670.120 ;
        RECT 4.400 636.800 1196.000 638.200 ;
        RECT 4.000 592.640 1196.000 636.800 ;
        RECT 4.000 591.240 1195.600 592.640 ;
        RECT 4.000 563.400 1196.000 591.240 ;
        RECT 4.400 562.000 1196.000 563.400 ;
        RECT 4.000 513.760 1196.000 562.000 ;
        RECT 4.000 512.360 1195.600 513.760 ;
        RECT 4.000 487.920 1196.000 512.360 ;
        RECT 4.400 486.520 1196.000 487.920 ;
        RECT 4.000 434.880 1196.000 486.520 ;
        RECT 4.000 433.480 1195.600 434.880 ;
        RECT 4.000 413.120 1196.000 433.480 ;
        RECT 4.400 411.720 1196.000 413.120 ;
        RECT 4.000 356.000 1196.000 411.720 ;
        RECT 4.000 354.600 1195.600 356.000 ;
        RECT 4.000 338.320 1196.000 354.600 ;
        RECT 4.400 336.920 1196.000 338.320 ;
        RECT 4.000 277.120 1196.000 336.920 ;
        RECT 4.000 275.720 1195.600 277.120 ;
        RECT 4.000 262.840 1196.000 275.720 ;
        RECT 4.400 261.440 1196.000 262.840 ;
        RECT 4.000 198.240 1196.000 261.440 ;
        RECT 4.000 196.840 1195.600 198.240 ;
        RECT 4.000 188.040 1196.000 196.840 ;
        RECT 4.400 186.640 1196.000 188.040 ;
        RECT 4.000 119.360 1196.000 186.640 ;
        RECT 4.000 117.960 1195.600 119.360 ;
        RECT 4.000 113.240 1196.000 117.960 ;
        RECT 4.400 111.840 1196.000 113.240 ;
        RECT 4.000 40.480 1196.000 111.840 ;
        RECT 4.000 39.080 1195.600 40.480 ;
        RECT 4.000 38.440 1196.000 39.080 ;
        RECT 4.400 37.040 1196.000 38.440 ;
        RECT 4.000 10.715 1196.000 37.040 ;
      LAYER met4 ;
        RECT 96.895 59.335 97.440 1484.265 ;
        RECT 99.840 59.335 174.240 1484.265 ;
        RECT 176.640 59.335 251.040 1484.265 ;
        RECT 253.440 59.335 327.840 1484.265 ;
        RECT 330.240 59.335 404.640 1484.265 ;
        RECT 407.040 59.335 481.440 1484.265 ;
        RECT 483.840 59.335 558.240 1484.265 ;
        RECT 560.640 59.335 635.040 1484.265 ;
        RECT 637.440 59.335 711.840 1484.265 ;
        RECT 714.240 59.335 788.640 1484.265 ;
        RECT 791.040 59.335 865.440 1484.265 ;
        RECT 867.840 59.335 942.240 1484.265 ;
        RECT 944.640 59.335 1019.040 1484.265 ;
        RECT 1021.440 59.335 1095.840 1484.265 ;
        RECT 1098.240 59.335 1132.225 1484.265 ;
  END
END custom_sram
END LIBRARY

