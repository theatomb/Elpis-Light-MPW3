VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO io_input_arbiter
  CLASS BLOCK ;
  FOREIGN io_input_arbiter ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 75.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END clk
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 71.000 30.730 75.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 71.000 35.330 75.000 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 71.000 54.190 75.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 40.840 75.000 41.440 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 71.000 63.390 75.000 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 63.280 75.000 63.880 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 71.000 67.990 75.000 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 71.000 11.870 75.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 71.000 16.470 75.000 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 25.880 75.000 26.480 ;
    END
  END data_out[9]
  PIN is_ready_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 71.000 2.670 75.000 ;
    END
  END is_ready_core0
  PIN read_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END read_enable
  PIN read_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 71.000 7.270 75.000 ;
    END
  END read_value[0]
  PIN read_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END read_value[10]
  PIN read_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END read_value[11]
  PIN read_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END read_value[12]
  PIN read_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END read_value[13]
  PIN read_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 33.360 75.000 33.960 ;
    END
  END read_value[14]
  PIN read_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 71.000 39.930 75.000 ;
    END
  END read_value[15]
  PIN read_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END read_value[16]
  PIN read_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 71.000 44.530 75.000 ;
    END
  END read_value[17]
  PIN read_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 71.000 49.130 75.000 ;
    END
  END read_value[18]
  PIN read_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END read_value[19]
  PIN read_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END read_value[1]
  PIN read_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END read_value[20]
  PIN read_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END read_value[21]
  PIN read_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END read_value[22]
  PIN read_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END read_value[23]
  PIN read_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 71.000 58.790 75.000 ;
    END
  END read_value[24]
  PIN read_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END read_value[25]
  PIN read_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 48.320 75.000 48.920 ;
    END
  END read_value[26]
  PIN read_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 55.800 75.000 56.400 ;
    END
  END read_value[27]
  PIN read_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 70.760 75.000 71.360 ;
    END
  END read_value[28]
  PIN read_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END read_value[29]
  PIN read_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END read_value[2]
  PIN read_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END read_value[30]
  PIN read_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 71.000 72.590 75.000 ;
    END
  END read_value[31]
  PIN read_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END read_value[3]
  PIN read_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 3.440 75.000 4.040 ;
    END
  END read_value[4]
  PIN read_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END read_value[5]
  PIN read_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 10.920 75.000 11.520 ;
    END
  END read_value[6]
  PIN read_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 71.000 21.070 75.000 ;
    END
  END read_value[7]
  PIN read_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 18.400 75.000 19.000 ;
    END
  END read_value[8]
  PIN read_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 71.000 25.670 75.000 ;
    END
  END read_value[9]
  PIN req_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END req_core0
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.380 10.640 16.980 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.700 10.640 38.300 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.020 10.640 59.620 62.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.040 10.640 27.640 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.360 10.640 48.960 62.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 3.825 70.695 62.645 ;
      LAYER met1 ;
        RECT 1.910 3.780 73.070 62.800 ;
      LAYER met2 ;
        RECT 1.940 70.720 2.110 73.285 ;
        RECT 2.950 70.720 6.710 73.285 ;
        RECT 7.550 70.720 11.310 73.285 ;
        RECT 12.150 70.720 15.910 73.285 ;
        RECT 16.750 70.720 20.510 73.285 ;
        RECT 21.350 70.720 25.110 73.285 ;
        RECT 25.950 70.720 30.170 73.285 ;
        RECT 31.010 70.720 34.770 73.285 ;
        RECT 35.610 70.720 39.370 73.285 ;
        RECT 40.210 70.720 43.970 73.285 ;
        RECT 44.810 70.720 48.570 73.285 ;
        RECT 49.410 70.720 53.630 73.285 ;
        RECT 54.470 70.720 58.230 73.285 ;
        RECT 59.070 70.720 62.830 73.285 ;
        RECT 63.670 70.720 67.430 73.285 ;
        RECT 68.270 70.720 72.030 73.285 ;
        RECT 72.870 70.720 73.040 73.285 ;
        RECT 1.940 4.280 73.040 70.720 ;
        RECT 2.490 1.515 5.330 4.280 ;
        RECT 6.170 1.515 9.010 4.280 ;
        RECT 9.850 1.515 12.690 4.280 ;
        RECT 13.530 1.515 16.370 4.280 ;
        RECT 17.210 1.515 20.050 4.280 ;
        RECT 20.890 1.515 23.730 4.280 ;
        RECT 24.570 1.515 27.870 4.280 ;
        RECT 28.710 1.515 31.550 4.280 ;
        RECT 32.390 1.515 35.230 4.280 ;
        RECT 36.070 1.515 38.910 4.280 ;
        RECT 39.750 1.515 42.590 4.280 ;
        RECT 43.430 1.515 46.270 4.280 ;
        RECT 47.110 1.515 49.950 4.280 ;
        RECT 50.790 1.515 54.090 4.280 ;
        RECT 54.930 1.515 57.770 4.280 ;
        RECT 58.610 1.515 61.450 4.280 ;
        RECT 62.290 1.515 65.130 4.280 ;
        RECT 65.970 1.515 68.810 4.280 ;
        RECT 69.650 1.515 72.490 4.280 ;
      LAYER met3 ;
        RECT 4.400 72.400 71.000 73.265 ;
        RECT 4.000 71.760 71.000 72.400 ;
        RECT 4.000 70.400 70.600 71.760 ;
        RECT 4.400 70.360 70.600 70.400 ;
        RECT 4.400 69.000 71.000 70.360 ;
        RECT 4.000 67.000 71.000 69.000 ;
        RECT 4.400 65.600 71.000 67.000 ;
        RECT 4.000 64.280 71.000 65.600 ;
        RECT 4.000 63.600 70.600 64.280 ;
        RECT 4.400 62.880 70.600 63.600 ;
        RECT 4.400 62.200 71.000 62.880 ;
        RECT 4.000 60.880 71.000 62.200 ;
        RECT 4.400 59.480 71.000 60.880 ;
        RECT 4.000 57.480 71.000 59.480 ;
        RECT 4.400 56.800 71.000 57.480 ;
        RECT 4.400 56.080 70.600 56.800 ;
        RECT 4.000 55.400 70.600 56.080 ;
        RECT 4.000 54.080 71.000 55.400 ;
        RECT 4.400 52.680 71.000 54.080 ;
        RECT 4.000 50.680 71.000 52.680 ;
        RECT 4.400 49.320 71.000 50.680 ;
        RECT 4.400 49.280 70.600 49.320 ;
        RECT 4.000 47.920 70.600 49.280 ;
        RECT 4.000 47.280 71.000 47.920 ;
        RECT 4.400 45.880 71.000 47.280 ;
        RECT 4.000 44.560 71.000 45.880 ;
        RECT 4.400 43.160 71.000 44.560 ;
        RECT 4.000 41.840 71.000 43.160 ;
        RECT 4.000 41.160 70.600 41.840 ;
        RECT 4.400 40.440 70.600 41.160 ;
        RECT 4.400 39.760 71.000 40.440 ;
        RECT 4.000 37.760 71.000 39.760 ;
        RECT 4.400 36.360 71.000 37.760 ;
        RECT 4.000 34.360 71.000 36.360 ;
        RECT 4.400 32.960 70.600 34.360 ;
        RECT 4.000 31.640 71.000 32.960 ;
        RECT 4.400 30.240 71.000 31.640 ;
        RECT 4.000 28.240 71.000 30.240 ;
        RECT 4.400 26.880 71.000 28.240 ;
        RECT 4.400 26.840 70.600 26.880 ;
        RECT 4.000 25.480 70.600 26.840 ;
        RECT 4.000 24.840 71.000 25.480 ;
        RECT 4.400 23.440 71.000 24.840 ;
        RECT 4.000 21.440 71.000 23.440 ;
        RECT 4.400 20.040 71.000 21.440 ;
        RECT 4.000 19.400 71.000 20.040 ;
        RECT 4.000 18.040 70.600 19.400 ;
        RECT 4.400 18.000 70.600 18.040 ;
        RECT 4.400 16.640 71.000 18.000 ;
        RECT 4.000 15.320 71.000 16.640 ;
        RECT 4.400 13.920 71.000 15.320 ;
        RECT 4.000 11.920 71.000 13.920 ;
        RECT 4.400 10.520 70.600 11.920 ;
        RECT 4.000 8.520 71.000 10.520 ;
        RECT 4.400 7.120 71.000 8.520 ;
        RECT 4.000 5.120 71.000 7.120 ;
        RECT 4.400 4.440 71.000 5.120 ;
        RECT 4.400 3.720 70.600 4.440 ;
        RECT 4.000 3.040 70.600 3.720 ;
        RECT 4.000 2.400 71.000 3.040 ;
        RECT 4.400 1.535 71.000 2.400 ;
  END
END io_input_arbiter
END LIBRARY

