VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.800 4.000 1195.400 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1215.880 1500.000 1216.480 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 0.000 1316.430 4.000 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 0.000 1333.910 4.000 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1277.080 4.000 1277.680 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1252.600 1500.000 1253.200 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1310.400 4.000 1311.000 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.720 4.000 1327.320 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.550 0.000 1403.830 4.000 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 0.000 1421.310 4.000 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.950 1496.000 1376.230 1500.000 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1359.360 4.000 1359.960 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.510 1496.000 1392.790 1500.000 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.510 0.000 1438.790 4.000 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.470 0.000 1473.750 4.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1343.720 1500.000 1344.320 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1362.080 1500.000 1362.680 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.170 1496.000 1425.450 1500.000 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 155.080 1500.000 155.680 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1380.440 1500.000 1381.040 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1442.320 4.000 1442.920 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.290 1496.000 1458.570 1500.000 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 1496.000 1475.130 1500.000 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1398.800 1500.000 1399.400 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1417.160 1500.000 1417.760 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1435.520 1500.000 1436.120 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1472.240 1500.000 1472.840 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 1496.000 403.790 1500.000 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 1496.000 453.010 1500.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 1496.000 502.690 1500.000 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 301.280 1500.000 301.880 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 1496.000 551.910 1500.000 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 392.400 1500.000 393.000 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 429.120 1500.000 429.720 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 465.840 1500.000 466.440 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 1496.000 601.590 1500.000 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 484.200 1500.000 484.800 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 1496.000 700.490 1500.000 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 557.640 1500.000 558.240 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 1496.000 766.270 1500.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 1496.000 782.830 1500.000 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 612.040 1500.000 612.640 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 0.000 793.410 4.000 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 634.480 4.000 635.080 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 667.120 1500.000 667.720 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 685.480 1500.000 686.080 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.120 4.000 667.720 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 4.000 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 1496.000 832.050 1500.000 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 740.560 1500.000 741.160 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.070 0.000 880.350 4.000 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 1496.000 898.290 1500.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 1496.000 172.870 1500.000 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.110 1496.000 914.390 1500.000 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 0.000 932.790 4.000 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 1496.000 930.950 1500.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 794.960 1500.000 795.560 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 766.400 4.000 767.000 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 4.000 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 1496.000 964.070 1500.000 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 1496.000 222.090 1500.000 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 1496.000 997.190 1500.000 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 1496.000 1013.290 1500.000 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 868.400 1500.000 869.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 886.760 1500.000 887.360 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.870 0.000 1055.150 4.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 1496.000 1062.970 1500.000 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 100.000 1500.000 100.600 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 905.120 1500.000 905.720 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 0.000 1124.610 4.000 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 923.480 1500.000 924.080 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.280 4.000 947.880 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 941.840 1500.000 942.440 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 1496.000 1128.750 1500.000 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 1496.000 1145.310 1500.000 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 996.240 1500.000 996.840 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.590 1496.000 1161.870 1500.000 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.150 1496.000 1178.430 1500.000 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1051.320 1500.000 1051.920 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1088.040 1500.000 1088.640 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 1496.000 1194.990 1500.000 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1124.760 1500.000 1125.360 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.730 0.000 1212.010 4.000 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1095.520 4.000 1096.120 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.930 1496.000 1244.210 1500.000 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1112.520 4.000 1113.120 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.160 4.000 1145.760 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 0.000 1246.970 4.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1160.800 1500.000 1161.400 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1161.480 4.000 1162.080 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.610 1496.000 1293.890 1500.000 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1178.480 4.000 1179.080 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 0.000 1281.930 4.000 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.670 0.000 1298.950 4.000 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1496.000 90.530 1500.000 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 1496.000 354.110 1500.000 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 1496.000 419.890 1500.000 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 246.200 1500.000 246.800 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 1496.000 486.130 1500.000 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 264.560 1500.000 265.160 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 26.560 1500.000 27.160 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 447.480 1500.000 448.080 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 1496.000 568.470 1500.000 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 1496.000 617.690 1500.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 1496.000 667.370 1500.000 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 502.560 1500.000 503.160 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 551.520 4.000 552.120 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 1496.000 123.190 1500.000 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 575.320 1500.000 575.920 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 1496.000 238.650 1500.000 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 1496.000 320.990 1500.000 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 1496.000 40.850 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 1496.000 73.970 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 1496.000 57.410 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 1496.000 337.550 1500.000 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 1496.000 370.670 1500.000 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 209.480 1500.000 210.080 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 1496.000 518.790 1500.000 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 319.640 1500.000 320.240 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 44.920 1500.000 45.520 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 63.280 1500.000 63.880 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 1496.000 271.770 1500.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 1496.000 107.090 1500.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1211.120 4.000 1211.720 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1244.440 4.000 1245.040 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1260.760 4.000 1261.360 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 1496.000 1343.110 1500.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.110 0.000 1351.390 4.000 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1234.240 1500.000 1234.840 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.390 1496.000 1359.670 1500.000 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.070 0.000 1386.350 4.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1270.960 1500.000 1271.560 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1289.320 1500.000 1289.920 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1307.680 1500.000 1308.280 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1376.360 4.000 1376.960 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.610 1496.000 1408.890 1500.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 0.000 1456.270 4.000 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1325.360 1500.000 1325.960 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.680 4.000 1393.280 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.000 4.000 1409.600 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 173.440 1500.000 174.040 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1425.320 4.000 1425.920 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.730 1496.000 1442.010 1500.000 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 1496.000 1491.690 1500.000 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1474.960 4.000 1475.560 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.280 4.000 1491.880 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1453.880 1500.000 1454.480 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1490.600 1500.000 1491.200 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 1496.000 436.450 1500.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 338.000 1500.000 338.600 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 356.360 1500.000 356.960 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 410.760 1500.000 411.360 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 1496.000 650.810 1500.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 1496.000 683.930 1500.000 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 1496.000 716.590 1500.000 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 539.280 1500.000 539.880 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 1496.000 139.750 1500.000 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 1496.000 749.710 1500.000 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 630.400 1500.000 631.000 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 1496.000 799.390 1500.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 648.760 1500.000 649.360 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 4.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 1496.000 815.490 1500.000 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 703.840 1500.000 704.440 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 722.200 1500.000 722.800 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 1496.000 848.610 1500.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 1496.000 865.170 1500.000 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 1496.000 881.730 1500.000 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 0.000 915.310 4.000 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 1496.000 189.430 1500.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 758.920 1500.000 759.520 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 4.000 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 776.600 1500.000 777.200 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 1496.000 947.510 1500.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 813.320 1500.000 813.920 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 1496.000 980.630 1500.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 0.000 1020.190 4.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 831.680 1500.000 832.280 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 1496.000 1029.850 1500.000 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 850.040 1500.000 850.640 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 1496.000 1046.410 1500.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 898.320 4.000 898.920 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 0.000 1089.650 4.000 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 0.000 1107.130 4.000 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 1496.000 1079.530 1500.000 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 1496.000 1096.090 1500.000 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.810 0.000 1142.090 4.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 1496.000 1112.190 1500.000 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.280 4.000 964.880 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 959.520 1500.000 960.120 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 4.000 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 977.880 1500.000 978.480 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 1496.000 288.330 1500.000 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1014.600 1500.000 1015.200 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1032.960 1500.000 1033.560 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1046.560 4.000 1047.160 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.880 4.000 1063.480 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1069.680 1500.000 1070.280 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1106.400 1500.000 1107.000 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1079.200 4.000 1079.800 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 1496.000 1211.090 1500.000 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 1496.000 1227.650 1500.000 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 118.360 1500.000 118.960 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.210 0.000 1229.490 4.000 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1142.440 1500.000 1143.040 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.490 1496.000 1260.770 1500.000 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 0.000 1264.450 4.000 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.050 1496.000 1277.330 1500.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 1496.000 1309.990 1500.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1179.160 1500.000 1179.760 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.270 1496.000 1326.550 1500.000 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1197.520 1500.000 1198.120 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 1496.000 8.190 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 1496.000 24.290 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 8.880 1500.000 9.480 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 191.800 1500.000 192.400 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 1496.000 387.230 1500.000 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 227.840 1500.000 228.440 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 1496.000 469.570 1500.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 282.920 1500.000 283.520 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 1496.000 535.350 1500.000 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 374.720 1500.000 375.320 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 1496.000 585.030 1500.000 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 1496.000 634.250 1500.000 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 1496.000 733.150 1500.000 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 520.920 1500.000 521.520 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 1496.000 156.310 1500.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 593.680 1500.000 594.280 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 1496.000 205.990 1500.000 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 81.640 1500.000 82.240 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 1496.000 255.210 1500.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 1496.000 304.890 1500.000 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 136.720 1500.000 137.320 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 7.520 1494.080 1489.160 ;
      LAYER met2 ;
        RECT 6.990 1495.720 7.630 1496.410 ;
        RECT 8.470 1495.720 23.730 1496.410 ;
        RECT 24.570 1495.720 40.290 1496.410 ;
        RECT 41.130 1495.720 56.850 1496.410 ;
        RECT 57.690 1495.720 73.410 1496.410 ;
        RECT 74.250 1495.720 89.970 1496.410 ;
        RECT 90.810 1495.720 106.530 1496.410 ;
        RECT 107.370 1495.720 122.630 1496.410 ;
        RECT 123.470 1495.720 139.190 1496.410 ;
        RECT 140.030 1495.720 155.750 1496.410 ;
        RECT 156.590 1495.720 172.310 1496.410 ;
        RECT 173.150 1495.720 188.870 1496.410 ;
        RECT 189.710 1495.720 205.430 1496.410 ;
        RECT 206.270 1495.720 221.530 1496.410 ;
        RECT 222.370 1495.720 238.090 1496.410 ;
        RECT 238.930 1495.720 254.650 1496.410 ;
        RECT 255.490 1495.720 271.210 1496.410 ;
        RECT 272.050 1495.720 287.770 1496.410 ;
        RECT 288.610 1495.720 304.330 1496.410 ;
        RECT 305.170 1495.720 320.430 1496.410 ;
        RECT 321.270 1495.720 336.990 1496.410 ;
        RECT 337.830 1495.720 353.550 1496.410 ;
        RECT 354.390 1495.720 370.110 1496.410 ;
        RECT 370.950 1495.720 386.670 1496.410 ;
        RECT 387.510 1495.720 403.230 1496.410 ;
        RECT 404.070 1495.720 419.330 1496.410 ;
        RECT 420.170 1495.720 435.890 1496.410 ;
        RECT 436.730 1495.720 452.450 1496.410 ;
        RECT 453.290 1495.720 469.010 1496.410 ;
        RECT 469.850 1495.720 485.570 1496.410 ;
        RECT 486.410 1495.720 502.130 1496.410 ;
        RECT 502.970 1495.720 518.230 1496.410 ;
        RECT 519.070 1495.720 534.790 1496.410 ;
        RECT 535.630 1495.720 551.350 1496.410 ;
        RECT 552.190 1495.720 567.910 1496.410 ;
        RECT 568.750 1495.720 584.470 1496.410 ;
        RECT 585.310 1495.720 601.030 1496.410 ;
        RECT 601.870 1495.720 617.130 1496.410 ;
        RECT 617.970 1495.720 633.690 1496.410 ;
        RECT 634.530 1495.720 650.250 1496.410 ;
        RECT 651.090 1495.720 666.810 1496.410 ;
        RECT 667.650 1495.720 683.370 1496.410 ;
        RECT 684.210 1495.720 699.930 1496.410 ;
        RECT 700.770 1495.720 716.030 1496.410 ;
        RECT 716.870 1495.720 732.590 1496.410 ;
        RECT 733.430 1495.720 749.150 1496.410 ;
        RECT 749.990 1495.720 765.710 1496.410 ;
        RECT 766.550 1495.720 782.270 1496.410 ;
        RECT 783.110 1495.720 798.830 1496.410 ;
        RECT 799.670 1495.720 814.930 1496.410 ;
        RECT 815.770 1495.720 831.490 1496.410 ;
        RECT 832.330 1495.720 848.050 1496.410 ;
        RECT 848.890 1495.720 864.610 1496.410 ;
        RECT 865.450 1495.720 881.170 1496.410 ;
        RECT 882.010 1495.720 897.730 1496.410 ;
        RECT 898.570 1495.720 913.830 1496.410 ;
        RECT 914.670 1495.720 930.390 1496.410 ;
        RECT 931.230 1495.720 946.950 1496.410 ;
        RECT 947.790 1495.720 963.510 1496.410 ;
        RECT 964.350 1495.720 980.070 1496.410 ;
        RECT 980.910 1495.720 996.630 1496.410 ;
        RECT 997.470 1495.720 1012.730 1496.410 ;
        RECT 1013.570 1495.720 1029.290 1496.410 ;
        RECT 1030.130 1495.720 1045.850 1496.410 ;
        RECT 1046.690 1495.720 1062.410 1496.410 ;
        RECT 1063.250 1495.720 1078.970 1496.410 ;
        RECT 1079.810 1495.720 1095.530 1496.410 ;
        RECT 1096.370 1495.720 1111.630 1496.410 ;
        RECT 1112.470 1495.720 1128.190 1496.410 ;
        RECT 1129.030 1495.720 1144.750 1496.410 ;
        RECT 1145.590 1495.720 1161.310 1496.410 ;
        RECT 1162.150 1495.720 1177.870 1496.410 ;
        RECT 1178.710 1495.720 1194.430 1496.410 ;
        RECT 1195.270 1495.720 1210.530 1496.410 ;
        RECT 1211.370 1495.720 1227.090 1496.410 ;
        RECT 1227.930 1495.720 1243.650 1496.410 ;
        RECT 1244.490 1495.720 1260.210 1496.410 ;
        RECT 1261.050 1495.720 1276.770 1496.410 ;
        RECT 1277.610 1495.720 1293.330 1496.410 ;
        RECT 1294.170 1495.720 1309.430 1496.410 ;
        RECT 1310.270 1495.720 1325.990 1496.410 ;
        RECT 1326.830 1495.720 1342.550 1496.410 ;
        RECT 1343.390 1495.720 1359.110 1496.410 ;
        RECT 1359.950 1495.720 1375.670 1496.410 ;
        RECT 1376.510 1495.720 1392.230 1496.410 ;
        RECT 1393.070 1495.720 1408.330 1496.410 ;
        RECT 1409.170 1495.720 1424.890 1496.410 ;
        RECT 1425.730 1495.720 1441.450 1496.410 ;
        RECT 1442.290 1495.720 1458.010 1496.410 ;
        RECT 1458.850 1495.720 1474.570 1496.410 ;
        RECT 1475.410 1495.720 1491.130 1496.410 ;
        RECT 6.990 4.280 1491.680 1495.720 ;
        RECT 6.990 3.670 8.090 4.280 ;
        RECT 8.930 3.670 25.110 4.280 ;
        RECT 25.950 3.670 42.590 4.280 ;
        RECT 43.430 3.670 60.070 4.280 ;
        RECT 60.910 3.670 77.550 4.280 ;
        RECT 78.390 3.670 95.030 4.280 ;
        RECT 95.870 3.670 112.510 4.280 ;
        RECT 113.350 3.670 129.990 4.280 ;
        RECT 130.830 3.670 147.470 4.280 ;
        RECT 148.310 3.670 164.950 4.280 ;
        RECT 165.790 3.670 182.430 4.280 ;
        RECT 183.270 3.670 199.910 4.280 ;
        RECT 200.750 3.670 217.390 4.280 ;
        RECT 218.230 3.670 234.410 4.280 ;
        RECT 235.250 3.670 251.890 4.280 ;
        RECT 252.730 3.670 269.370 4.280 ;
        RECT 270.210 3.670 286.850 4.280 ;
        RECT 287.690 3.670 304.330 4.280 ;
        RECT 305.170 3.670 321.810 4.280 ;
        RECT 322.650 3.670 339.290 4.280 ;
        RECT 340.130 3.670 356.770 4.280 ;
        RECT 357.610 3.670 374.250 4.280 ;
        RECT 375.090 3.670 391.730 4.280 ;
        RECT 392.570 3.670 409.210 4.280 ;
        RECT 410.050 3.670 426.690 4.280 ;
        RECT 427.530 3.670 443.710 4.280 ;
        RECT 444.550 3.670 461.190 4.280 ;
        RECT 462.030 3.670 478.670 4.280 ;
        RECT 479.510 3.670 496.150 4.280 ;
        RECT 496.990 3.670 513.630 4.280 ;
        RECT 514.470 3.670 531.110 4.280 ;
        RECT 531.950 3.670 548.590 4.280 ;
        RECT 549.430 3.670 566.070 4.280 ;
        RECT 566.910 3.670 583.550 4.280 ;
        RECT 584.390 3.670 601.030 4.280 ;
        RECT 601.870 3.670 618.510 4.280 ;
        RECT 619.350 3.670 635.990 4.280 ;
        RECT 636.830 3.670 653.010 4.280 ;
        RECT 653.850 3.670 670.490 4.280 ;
        RECT 671.330 3.670 687.970 4.280 ;
        RECT 688.810 3.670 705.450 4.280 ;
        RECT 706.290 3.670 722.930 4.280 ;
        RECT 723.770 3.670 740.410 4.280 ;
        RECT 741.250 3.670 757.890 4.280 ;
        RECT 758.730 3.670 775.370 4.280 ;
        RECT 776.210 3.670 792.850 4.280 ;
        RECT 793.690 3.670 810.330 4.280 ;
        RECT 811.170 3.670 827.810 4.280 ;
        RECT 828.650 3.670 845.290 4.280 ;
        RECT 846.130 3.670 862.770 4.280 ;
        RECT 863.610 3.670 879.790 4.280 ;
        RECT 880.630 3.670 897.270 4.280 ;
        RECT 898.110 3.670 914.750 4.280 ;
        RECT 915.590 3.670 932.230 4.280 ;
        RECT 933.070 3.670 949.710 4.280 ;
        RECT 950.550 3.670 967.190 4.280 ;
        RECT 968.030 3.670 984.670 4.280 ;
        RECT 985.510 3.670 1002.150 4.280 ;
        RECT 1002.990 3.670 1019.630 4.280 ;
        RECT 1020.470 3.670 1037.110 4.280 ;
        RECT 1037.950 3.670 1054.590 4.280 ;
        RECT 1055.430 3.670 1072.070 4.280 ;
        RECT 1072.910 3.670 1089.090 4.280 ;
        RECT 1089.930 3.670 1106.570 4.280 ;
        RECT 1107.410 3.670 1124.050 4.280 ;
        RECT 1124.890 3.670 1141.530 4.280 ;
        RECT 1142.370 3.670 1159.010 4.280 ;
        RECT 1159.850 3.670 1176.490 4.280 ;
        RECT 1177.330 3.670 1193.970 4.280 ;
        RECT 1194.810 3.670 1211.450 4.280 ;
        RECT 1212.290 3.670 1228.930 4.280 ;
        RECT 1229.770 3.670 1246.410 4.280 ;
        RECT 1247.250 3.670 1263.890 4.280 ;
        RECT 1264.730 3.670 1281.370 4.280 ;
        RECT 1282.210 3.670 1298.390 4.280 ;
        RECT 1299.230 3.670 1315.870 4.280 ;
        RECT 1316.710 3.670 1333.350 4.280 ;
        RECT 1334.190 3.670 1350.830 4.280 ;
        RECT 1351.670 3.670 1368.310 4.280 ;
        RECT 1369.150 3.670 1385.790 4.280 ;
        RECT 1386.630 3.670 1403.270 4.280 ;
        RECT 1404.110 3.670 1420.750 4.280 ;
        RECT 1421.590 3.670 1438.230 4.280 ;
        RECT 1439.070 3.670 1455.710 4.280 ;
        RECT 1456.550 3.670 1473.190 4.280 ;
        RECT 1474.030 3.670 1490.670 4.280 ;
        RECT 1491.510 3.670 1491.680 4.280 ;
      LAYER met3 ;
        RECT 4.400 1491.600 1496.000 1491.745 ;
        RECT 4.400 1490.880 1495.600 1491.600 ;
        RECT 4.000 1490.200 1495.600 1490.880 ;
        RECT 4.000 1475.960 1496.000 1490.200 ;
        RECT 4.400 1474.560 1496.000 1475.960 ;
        RECT 4.000 1473.240 1496.000 1474.560 ;
        RECT 4.000 1471.840 1495.600 1473.240 ;
        RECT 4.000 1459.640 1496.000 1471.840 ;
        RECT 4.400 1458.240 1496.000 1459.640 ;
        RECT 4.000 1454.880 1496.000 1458.240 ;
        RECT 4.000 1453.480 1495.600 1454.880 ;
        RECT 4.000 1443.320 1496.000 1453.480 ;
        RECT 4.400 1441.920 1496.000 1443.320 ;
        RECT 4.000 1436.520 1496.000 1441.920 ;
        RECT 4.000 1435.120 1495.600 1436.520 ;
        RECT 4.000 1426.320 1496.000 1435.120 ;
        RECT 4.400 1424.920 1496.000 1426.320 ;
        RECT 4.000 1418.160 1496.000 1424.920 ;
        RECT 4.000 1416.760 1495.600 1418.160 ;
        RECT 4.000 1410.000 1496.000 1416.760 ;
        RECT 4.400 1408.600 1496.000 1410.000 ;
        RECT 4.000 1399.800 1496.000 1408.600 ;
        RECT 4.000 1398.400 1495.600 1399.800 ;
        RECT 4.000 1393.680 1496.000 1398.400 ;
        RECT 4.400 1392.280 1496.000 1393.680 ;
        RECT 4.000 1381.440 1496.000 1392.280 ;
        RECT 4.000 1380.040 1495.600 1381.440 ;
        RECT 4.000 1377.360 1496.000 1380.040 ;
        RECT 4.400 1375.960 1496.000 1377.360 ;
        RECT 4.000 1363.080 1496.000 1375.960 ;
        RECT 4.000 1361.680 1495.600 1363.080 ;
        RECT 4.000 1360.360 1496.000 1361.680 ;
        RECT 4.400 1358.960 1496.000 1360.360 ;
        RECT 4.000 1344.720 1496.000 1358.960 ;
        RECT 4.000 1344.040 1495.600 1344.720 ;
        RECT 4.400 1343.320 1495.600 1344.040 ;
        RECT 4.400 1342.640 1496.000 1343.320 ;
        RECT 4.000 1327.720 1496.000 1342.640 ;
        RECT 4.400 1326.360 1496.000 1327.720 ;
        RECT 4.400 1326.320 1495.600 1326.360 ;
        RECT 4.000 1324.960 1495.600 1326.320 ;
        RECT 4.000 1311.400 1496.000 1324.960 ;
        RECT 4.400 1310.000 1496.000 1311.400 ;
        RECT 4.000 1308.680 1496.000 1310.000 ;
        RECT 4.000 1307.280 1495.600 1308.680 ;
        RECT 4.000 1294.400 1496.000 1307.280 ;
        RECT 4.400 1293.000 1496.000 1294.400 ;
        RECT 4.000 1290.320 1496.000 1293.000 ;
        RECT 4.000 1288.920 1495.600 1290.320 ;
        RECT 4.000 1278.080 1496.000 1288.920 ;
        RECT 4.400 1276.680 1496.000 1278.080 ;
        RECT 4.000 1271.960 1496.000 1276.680 ;
        RECT 4.000 1270.560 1495.600 1271.960 ;
        RECT 4.000 1261.760 1496.000 1270.560 ;
        RECT 4.400 1260.360 1496.000 1261.760 ;
        RECT 4.000 1253.600 1496.000 1260.360 ;
        RECT 4.000 1252.200 1495.600 1253.600 ;
        RECT 4.000 1245.440 1496.000 1252.200 ;
        RECT 4.400 1244.040 1496.000 1245.440 ;
        RECT 4.000 1235.240 1496.000 1244.040 ;
        RECT 4.000 1233.840 1495.600 1235.240 ;
        RECT 4.000 1228.440 1496.000 1233.840 ;
        RECT 4.400 1227.040 1496.000 1228.440 ;
        RECT 4.000 1216.880 1496.000 1227.040 ;
        RECT 4.000 1215.480 1495.600 1216.880 ;
        RECT 4.000 1212.120 1496.000 1215.480 ;
        RECT 4.400 1210.720 1496.000 1212.120 ;
        RECT 4.000 1198.520 1496.000 1210.720 ;
        RECT 4.000 1197.120 1495.600 1198.520 ;
        RECT 4.000 1195.800 1496.000 1197.120 ;
        RECT 4.400 1194.400 1496.000 1195.800 ;
        RECT 4.000 1180.160 1496.000 1194.400 ;
        RECT 4.000 1179.480 1495.600 1180.160 ;
        RECT 4.400 1178.760 1495.600 1179.480 ;
        RECT 4.400 1178.080 1496.000 1178.760 ;
        RECT 4.000 1162.480 1496.000 1178.080 ;
        RECT 4.400 1161.800 1496.000 1162.480 ;
        RECT 4.400 1161.080 1495.600 1161.800 ;
        RECT 4.000 1160.400 1495.600 1161.080 ;
        RECT 4.000 1146.160 1496.000 1160.400 ;
        RECT 4.400 1144.760 1496.000 1146.160 ;
        RECT 4.000 1143.440 1496.000 1144.760 ;
        RECT 4.000 1142.040 1495.600 1143.440 ;
        RECT 4.000 1129.840 1496.000 1142.040 ;
        RECT 4.400 1128.440 1496.000 1129.840 ;
        RECT 4.000 1125.760 1496.000 1128.440 ;
        RECT 4.000 1124.360 1495.600 1125.760 ;
        RECT 4.000 1113.520 1496.000 1124.360 ;
        RECT 4.400 1112.120 1496.000 1113.520 ;
        RECT 4.000 1107.400 1496.000 1112.120 ;
        RECT 4.000 1106.000 1495.600 1107.400 ;
        RECT 4.000 1096.520 1496.000 1106.000 ;
        RECT 4.400 1095.120 1496.000 1096.520 ;
        RECT 4.000 1089.040 1496.000 1095.120 ;
        RECT 4.000 1087.640 1495.600 1089.040 ;
        RECT 4.000 1080.200 1496.000 1087.640 ;
        RECT 4.400 1078.800 1496.000 1080.200 ;
        RECT 4.000 1070.680 1496.000 1078.800 ;
        RECT 4.000 1069.280 1495.600 1070.680 ;
        RECT 4.000 1063.880 1496.000 1069.280 ;
        RECT 4.400 1062.480 1496.000 1063.880 ;
        RECT 4.000 1052.320 1496.000 1062.480 ;
        RECT 4.000 1050.920 1495.600 1052.320 ;
        RECT 4.000 1047.560 1496.000 1050.920 ;
        RECT 4.400 1046.160 1496.000 1047.560 ;
        RECT 4.000 1033.960 1496.000 1046.160 ;
        RECT 4.000 1032.560 1495.600 1033.960 ;
        RECT 4.000 1030.560 1496.000 1032.560 ;
        RECT 4.400 1029.160 1496.000 1030.560 ;
        RECT 4.000 1015.600 1496.000 1029.160 ;
        RECT 4.000 1014.240 1495.600 1015.600 ;
        RECT 4.400 1014.200 1495.600 1014.240 ;
        RECT 4.400 1012.840 1496.000 1014.200 ;
        RECT 4.000 997.920 1496.000 1012.840 ;
        RECT 4.400 997.240 1496.000 997.920 ;
        RECT 4.400 996.520 1495.600 997.240 ;
        RECT 4.000 995.840 1495.600 996.520 ;
        RECT 4.000 981.600 1496.000 995.840 ;
        RECT 4.400 980.200 1496.000 981.600 ;
        RECT 4.000 978.880 1496.000 980.200 ;
        RECT 4.000 977.480 1495.600 978.880 ;
        RECT 4.000 965.280 1496.000 977.480 ;
        RECT 4.400 963.880 1496.000 965.280 ;
        RECT 4.000 960.520 1496.000 963.880 ;
        RECT 4.000 959.120 1495.600 960.520 ;
        RECT 4.000 948.280 1496.000 959.120 ;
        RECT 4.400 946.880 1496.000 948.280 ;
        RECT 4.000 942.840 1496.000 946.880 ;
        RECT 4.000 941.440 1495.600 942.840 ;
        RECT 4.000 931.960 1496.000 941.440 ;
        RECT 4.400 930.560 1496.000 931.960 ;
        RECT 4.000 924.480 1496.000 930.560 ;
        RECT 4.000 923.080 1495.600 924.480 ;
        RECT 4.000 915.640 1496.000 923.080 ;
        RECT 4.400 914.240 1496.000 915.640 ;
        RECT 4.000 906.120 1496.000 914.240 ;
        RECT 4.000 904.720 1495.600 906.120 ;
        RECT 4.000 899.320 1496.000 904.720 ;
        RECT 4.400 897.920 1496.000 899.320 ;
        RECT 4.000 887.760 1496.000 897.920 ;
        RECT 4.000 886.360 1495.600 887.760 ;
        RECT 4.000 882.320 1496.000 886.360 ;
        RECT 4.400 880.920 1496.000 882.320 ;
        RECT 4.000 869.400 1496.000 880.920 ;
        RECT 4.000 868.000 1495.600 869.400 ;
        RECT 4.000 866.000 1496.000 868.000 ;
        RECT 4.400 864.600 1496.000 866.000 ;
        RECT 4.000 851.040 1496.000 864.600 ;
        RECT 4.000 849.680 1495.600 851.040 ;
        RECT 4.400 849.640 1495.600 849.680 ;
        RECT 4.400 848.280 1496.000 849.640 ;
        RECT 4.000 833.360 1496.000 848.280 ;
        RECT 4.400 832.680 1496.000 833.360 ;
        RECT 4.400 831.960 1495.600 832.680 ;
        RECT 4.000 831.280 1495.600 831.960 ;
        RECT 4.000 816.360 1496.000 831.280 ;
        RECT 4.400 814.960 1496.000 816.360 ;
        RECT 4.000 814.320 1496.000 814.960 ;
        RECT 4.000 812.920 1495.600 814.320 ;
        RECT 4.000 800.040 1496.000 812.920 ;
        RECT 4.400 798.640 1496.000 800.040 ;
        RECT 4.000 795.960 1496.000 798.640 ;
        RECT 4.000 794.560 1495.600 795.960 ;
        RECT 4.000 783.720 1496.000 794.560 ;
        RECT 4.400 782.320 1496.000 783.720 ;
        RECT 4.000 777.600 1496.000 782.320 ;
        RECT 4.000 776.200 1495.600 777.600 ;
        RECT 4.000 767.400 1496.000 776.200 ;
        RECT 4.400 766.000 1496.000 767.400 ;
        RECT 4.000 759.920 1496.000 766.000 ;
        RECT 4.000 758.520 1495.600 759.920 ;
        RECT 4.000 750.400 1496.000 758.520 ;
        RECT 4.400 749.000 1496.000 750.400 ;
        RECT 4.000 741.560 1496.000 749.000 ;
        RECT 4.000 740.160 1495.600 741.560 ;
        RECT 4.000 734.080 1496.000 740.160 ;
        RECT 4.400 732.680 1496.000 734.080 ;
        RECT 4.000 723.200 1496.000 732.680 ;
        RECT 4.000 721.800 1495.600 723.200 ;
        RECT 4.000 717.760 1496.000 721.800 ;
        RECT 4.400 716.360 1496.000 717.760 ;
        RECT 4.000 704.840 1496.000 716.360 ;
        RECT 4.000 703.440 1495.600 704.840 ;
        RECT 4.000 701.440 1496.000 703.440 ;
        RECT 4.400 700.040 1496.000 701.440 ;
        RECT 4.000 686.480 1496.000 700.040 ;
        RECT 4.000 685.080 1495.600 686.480 ;
        RECT 4.000 684.440 1496.000 685.080 ;
        RECT 4.400 683.040 1496.000 684.440 ;
        RECT 4.000 668.120 1496.000 683.040 ;
        RECT 4.400 666.720 1495.600 668.120 ;
        RECT 4.000 651.800 1496.000 666.720 ;
        RECT 4.400 650.400 1496.000 651.800 ;
        RECT 4.000 649.760 1496.000 650.400 ;
        RECT 4.000 648.360 1495.600 649.760 ;
        RECT 4.000 635.480 1496.000 648.360 ;
        RECT 4.400 634.080 1496.000 635.480 ;
        RECT 4.000 631.400 1496.000 634.080 ;
        RECT 4.000 630.000 1495.600 631.400 ;
        RECT 4.000 618.480 1496.000 630.000 ;
        RECT 4.400 617.080 1496.000 618.480 ;
        RECT 4.000 613.040 1496.000 617.080 ;
        RECT 4.000 611.640 1495.600 613.040 ;
        RECT 4.000 602.160 1496.000 611.640 ;
        RECT 4.400 600.760 1496.000 602.160 ;
        RECT 4.000 594.680 1496.000 600.760 ;
        RECT 4.000 593.280 1495.600 594.680 ;
        RECT 4.000 585.840 1496.000 593.280 ;
        RECT 4.400 584.440 1496.000 585.840 ;
        RECT 4.000 576.320 1496.000 584.440 ;
        RECT 4.000 574.920 1495.600 576.320 ;
        RECT 4.000 569.520 1496.000 574.920 ;
        RECT 4.400 568.120 1496.000 569.520 ;
        RECT 4.000 558.640 1496.000 568.120 ;
        RECT 4.000 557.240 1495.600 558.640 ;
        RECT 4.000 552.520 1496.000 557.240 ;
        RECT 4.400 551.120 1496.000 552.520 ;
        RECT 4.000 540.280 1496.000 551.120 ;
        RECT 4.000 538.880 1495.600 540.280 ;
        RECT 4.000 536.200 1496.000 538.880 ;
        RECT 4.400 534.800 1496.000 536.200 ;
        RECT 4.000 521.920 1496.000 534.800 ;
        RECT 4.000 520.520 1495.600 521.920 ;
        RECT 4.000 519.880 1496.000 520.520 ;
        RECT 4.400 518.480 1496.000 519.880 ;
        RECT 4.000 503.560 1496.000 518.480 ;
        RECT 4.400 502.160 1495.600 503.560 ;
        RECT 4.000 487.240 1496.000 502.160 ;
        RECT 4.400 485.840 1496.000 487.240 ;
        RECT 4.000 485.200 1496.000 485.840 ;
        RECT 4.000 483.800 1495.600 485.200 ;
        RECT 4.000 470.240 1496.000 483.800 ;
        RECT 4.400 468.840 1496.000 470.240 ;
        RECT 4.000 466.840 1496.000 468.840 ;
        RECT 4.000 465.440 1495.600 466.840 ;
        RECT 4.000 453.920 1496.000 465.440 ;
        RECT 4.400 452.520 1496.000 453.920 ;
        RECT 4.000 448.480 1496.000 452.520 ;
        RECT 4.000 447.080 1495.600 448.480 ;
        RECT 4.000 437.600 1496.000 447.080 ;
        RECT 4.400 436.200 1496.000 437.600 ;
        RECT 4.000 430.120 1496.000 436.200 ;
        RECT 4.000 428.720 1495.600 430.120 ;
        RECT 4.000 421.280 1496.000 428.720 ;
        RECT 4.400 419.880 1496.000 421.280 ;
        RECT 4.000 411.760 1496.000 419.880 ;
        RECT 4.000 410.360 1495.600 411.760 ;
        RECT 4.000 404.280 1496.000 410.360 ;
        RECT 4.400 402.880 1496.000 404.280 ;
        RECT 4.000 393.400 1496.000 402.880 ;
        RECT 4.000 392.000 1495.600 393.400 ;
        RECT 4.000 387.960 1496.000 392.000 ;
        RECT 4.400 386.560 1496.000 387.960 ;
        RECT 4.000 375.720 1496.000 386.560 ;
        RECT 4.000 374.320 1495.600 375.720 ;
        RECT 4.000 371.640 1496.000 374.320 ;
        RECT 4.400 370.240 1496.000 371.640 ;
        RECT 4.000 357.360 1496.000 370.240 ;
        RECT 4.000 355.960 1495.600 357.360 ;
        RECT 4.000 355.320 1496.000 355.960 ;
        RECT 4.400 353.920 1496.000 355.320 ;
        RECT 4.000 339.000 1496.000 353.920 ;
        RECT 4.000 338.320 1495.600 339.000 ;
        RECT 4.400 337.600 1495.600 338.320 ;
        RECT 4.400 336.920 1496.000 337.600 ;
        RECT 4.000 322.000 1496.000 336.920 ;
        RECT 4.400 320.640 1496.000 322.000 ;
        RECT 4.400 320.600 1495.600 320.640 ;
        RECT 4.000 319.240 1495.600 320.600 ;
        RECT 4.000 305.680 1496.000 319.240 ;
        RECT 4.400 304.280 1496.000 305.680 ;
        RECT 4.000 302.280 1496.000 304.280 ;
        RECT 4.000 300.880 1495.600 302.280 ;
        RECT 4.000 289.360 1496.000 300.880 ;
        RECT 4.400 287.960 1496.000 289.360 ;
        RECT 4.000 283.920 1496.000 287.960 ;
        RECT 4.000 282.520 1495.600 283.920 ;
        RECT 4.000 272.360 1496.000 282.520 ;
        RECT 4.400 270.960 1496.000 272.360 ;
        RECT 4.000 265.560 1496.000 270.960 ;
        RECT 4.000 264.160 1495.600 265.560 ;
        RECT 4.000 256.040 1496.000 264.160 ;
        RECT 4.400 254.640 1496.000 256.040 ;
        RECT 4.000 247.200 1496.000 254.640 ;
        RECT 4.000 245.800 1495.600 247.200 ;
        RECT 4.000 239.720 1496.000 245.800 ;
        RECT 4.400 238.320 1496.000 239.720 ;
        RECT 4.000 228.840 1496.000 238.320 ;
        RECT 4.000 227.440 1495.600 228.840 ;
        RECT 4.000 223.400 1496.000 227.440 ;
        RECT 4.400 222.000 1496.000 223.400 ;
        RECT 4.000 210.480 1496.000 222.000 ;
        RECT 4.000 209.080 1495.600 210.480 ;
        RECT 4.000 206.400 1496.000 209.080 ;
        RECT 4.400 205.000 1496.000 206.400 ;
        RECT 4.000 192.800 1496.000 205.000 ;
        RECT 4.000 191.400 1495.600 192.800 ;
        RECT 4.000 190.080 1496.000 191.400 ;
        RECT 4.400 188.680 1496.000 190.080 ;
        RECT 4.000 174.440 1496.000 188.680 ;
        RECT 4.000 173.760 1495.600 174.440 ;
        RECT 4.400 173.040 1495.600 173.760 ;
        RECT 4.400 172.360 1496.000 173.040 ;
        RECT 4.000 157.440 1496.000 172.360 ;
        RECT 4.400 156.080 1496.000 157.440 ;
        RECT 4.400 156.040 1495.600 156.080 ;
        RECT 4.000 154.680 1495.600 156.040 ;
        RECT 4.000 140.440 1496.000 154.680 ;
        RECT 4.400 139.040 1496.000 140.440 ;
        RECT 4.000 137.720 1496.000 139.040 ;
        RECT 4.000 136.320 1495.600 137.720 ;
        RECT 4.000 124.120 1496.000 136.320 ;
        RECT 4.400 122.720 1496.000 124.120 ;
        RECT 4.000 119.360 1496.000 122.720 ;
        RECT 4.000 117.960 1495.600 119.360 ;
        RECT 4.000 107.800 1496.000 117.960 ;
        RECT 4.400 106.400 1496.000 107.800 ;
        RECT 4.000 101.000 1496.000 106.400 ;
        RECT 4.000 99.600 1495.600 101.000 ;
        RECT 4.000 91.480 1496.000 99.600 ;
        RECT 4.400 90.080 1496.000 91.480 ;
        RECT 4.000 82.640 1496.000 90.080 ;
        RECT 4.000 81.240 1495.600 82.640 ;
        RECT 4.000 74.480 1496.000 81.240 ;
        RECT 4.400 73.080 1496.000 74.480 ;
        RECT 4.000 64.280 1496.000 73.080 ;
        RECT 4.000 62.880 1495.600 64.280 ;
        RECT 4.000 58.160 1496.000 62.880 ;
        RECT 4.400 56.760 1496.000 58.160 ;
        RECT 4.000 45.920 1496.000 56.760 ;
        RECT 4.000 44.520 1495.600 45.920 ;
        RECT 4.000 41.840 1496.000 44.520 ;
        RECT 4.400 40.440 1496.000 41.840 ;
        RECT 4.000 27.560 1496.000 40.440 ;
        RECT 4.000 26.160 1495.600 27.560 ;
        RECT 4.000 25.520 1496.000 26.160 ;
        RECT 4.400 24.120 1496.000 25.520 ;
        RECT 4.000 9.880 1496.000 24.120 ;
        RECT 4.000 9.200 1495.600 9.880 ;
        RECT 4.400 8.480 1495.600 9.200 ;
        RECT 4.400 8.335 1496.000 8.480 ;
      LAYER met4 ;
        RECT 164.975 11.735 174.240 1486.305 ;
        RECT 176.640 11.735 251.040 1486.305 ;
        RECT 253.440 11.735 327.840 1486.305 ;
        RECT 330.240 11.735 404.640 1486.305 ;
        RECT 407.040 11.735 481.440 1486.305 ;
        RECT 483.840 11.735 558.240 1486.305 ;
        RECT 560.640 11.735 635.040 1486.305 ;
        RECT 637.440 11.735 711.840 1486.305 ;
        RECT 714.240 11.735 788.640 1486.305 ;
        RECT 791.040 11.735 865.440 1486.305 ;
        RECT 867.840 11.735 942.240 1486.305 ;
        RECT 944.640 11.735 1019.040 1486.305 ;
        RECT 1021.440 11.735 1031.945 1486.305 ;
  END
END core
END LIBRARY

