* NGSPICE file created from chip_controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_8 abstract view
.subckt sky130_fd_sc_hd__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_4 abstract view
.subckt sky130_fd_sc_hd__fill_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt chip_controller addr0_to_sram[0] addr0_to_sram[10] addr0_to_sram[11] addr0_to_sram[12]
+ addr0_to_sram[13] addr0_to_sram[14] addr0_to_sram[15] addr0_to_sram[16] addr0_to_sram[17]
+ addr0_to_sram[18] addr0_to_sram[19] addr0_to_sram[1] addr0_to_sram[2] addr0_to_sram[3]
+ addr0_to_sram[4] addr0_to_sram[5] addr0_to_sram[6] addr0_to_sram[7] addr0_to_sram[8]
+ addr0_to_sram[9] addr_in[0] addr_in[10] addr_in[11] addr_in[12] addr_in[13] addr_in[14]
+ addr_in[15] addr_in[16] addr_in[17] addr_in[18] addr_in[19] addr_in[1] addr_in[2]
+ addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in[8] addr_in[9] addr_to_core_mem[0]
+ addr_to_core_mem[10] addr_to_core_mem[11] addr_to_core_mem[12] addr_to_core_mem[13]
+ addr_to_core_mem[14] addr_to_core_mem[15] addr_to_core_mem[16] addr_to_core_mem[17]
+ addr_to_core_mem[18] addr_to_core_mem[19] addr_to_core_mem[1] addr_to_core_mem[2]
+ addr_to_core_mem[3] addr_to_core_mem[4] addr_to_core_mem[5] addr_to_core_mem[6]
+ addr_to_core_mem[7] addr_to_core_mem[8] addr_to_core_mem[9] clk core0_data_print[0]
+ core0_data_print[10] core0_data_print[11] core0_data_print[12] core0_data_print[13]
+ core0_data_print[14] core0_data_print[15] core0_data_print[16] core0_data_print[17]
+ core0_data_print[18] core0_data_print[19] core0_data_print[1] core0_data_print[20]
+ core0_data_print[21] core0_data_print[22] core0_data_print[23] core0_data_print[24]
+ core0_data_print[25] core0_data_print[26] core0_data_print[27] core0_data_print[28]
+ core0_data_print[29] core0_data_print[2] core0_data_print[30] core0_data_print[31]
+ core0_data_print[3] core0_data_print[4] core0_data_print[5] core0_data_print[6]
+ core0_data_print[7] core0_data_print[8] core0_data_print[9] csb0_to_sram data_out_to_core[0]
+ data_out_to_core[10] data_out_to_core[11] data_out_to_core[12] data_out_to_core[13]
+ data_out_to_core[14] data_out_to_core[15] data_out_to_core[16] data_out_to_core[17]
+ data_out_to_core[18] data_out_to_core[19] data_out_to_core[1] data_out_to_core[20]
+ data_out_to_core[21] data_out_to_core[22] data_out_to_core[23] data_out_to_core[24]
+ data_out_to_core[25] data_out_to_core[26] data_out_to_core[27] data_out_to_core[28]
+ data_out_to_core[29] data_out_to_core[2] data_out_to_core[30] data_out_to_core[31]
+ data_out_to_core[3] data_out_to_core[4] data_out_to_core[5] data_out_to_core[6]
+ data_out_to_core[7] data_out_to_core[8] data_out_to_core[9] data_to_core_mem[0]
+ data_to_core_mem[10] data_to_core_mem[11] data_to_core_mem[12] data_to_core_mem[13]
+ data_to_core_mem[14] data_to_core_mem[15] data_to_core_mem[16] data_to_core_mem[17]
+ data_to_core_mem[18] data_to_core_mem[19] data_to_core_mem[1] data_to_core_mem[20]
+ data_to_core_mem[21] data_to_core_mem[22] data_to_core_mem[23] data_to_core_mem[24]
+ data_to_core_mem[25] data_to_core_mem[26] data_to_core_mem[27] data_to_core_mem[28]
+ data_to_core_mem[29] data_to_core_mem[2] data_to_core_mem[30] data_to_core_mem[31]
+ data_to_core_mem[3] data_to_core_mem[4] data_to_core_mem[5] data_to_core_mem[6]
+ data_to_core_mem[7] data_to_core_mem[8] data_to_core_mem[9] din0_to_sram[0] din0_to_sram[10]
+ din0_to_sram[11] din0_to_sram[12] din0_to_sram[13] din0_to_sram[14] din0_to_sram[15]
+ din0_to_sram[16] din0_to_sram[17] din0_to_sram[18] din0_to_sram[19] din0_to_sram[1]
+ din0_to_sram[20] din0_to_sram[21] din0_to_sram[22] din0_to_sram[23] din0_to_sram[24]
+ din0_to_sram[25] din0_to_sram[26] din0_to_sram[27] din0_to_sram[28] din0_to_sram[29]
+ din0_to_sram[2] din0_to_sram[30] din0_to_sram[31] din0_to_sram[3] din0_to_sram[4]
+ din0_to_sram[5] din0_to_sram[6] din0_to_sram[7] din0_to_sram[8] din0_to_sram[9]
+ dout0_to_sram[0] dout0_to_sram[10] dout0_to_sram[11] dout0_to_sram[12] dout0_to_sram[13]
+ dout0_to_sram[14] dout0_to_sram[15] dout0_to_sram[16] dout0_to_sram[17] dout0_to_sram[18]
+ dout0_to_sram[19] dout0_to_sram[1] dout0_to_sram[20] dout0_to_sram[21] dout0_to_sram[22]
+ dout0_to_sram[23] dout0_to_sram[24] dout0_to_sram[25] dout0_to_sram[26] dout0_to_sram[27]
+ dout0_to_sram[28] dout0_to_sram[29] dout0_to_sram[2] dout0_to_sram[30] dout0_to_sram[31]
+ dout0_to_sram[3] dout0_to_sram[4] dout0_to_sram[5] dout0_to_sram[6] dout0_to_sram[7]
+ dout0_to_sram[8] dout0_to_sram[9] is_loading_memory_into_core is_ready_dataout_core0
+ is_ready_print_core0 la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] rd_data_out[0] rd_data_out[100] rd_data_out[101]
+ rd_data_out[102] rd_data_out[103] rd_data_out[104] rd_data_out[105] rd_data_out[106]
+ rd_data_out[107] rd_data_out[108] rd_data_out[109] rd_data_out[10] rd_data_out[110]
+ rd_data_out[111] rd_data_out[112] rd_data_out[113] rd_data_out[114] rd_data_out[115]
+ rd_data_out[116] rd_data_out[117] rd_data_out[118] rd_data_out[119] rd_data_out[11]
+ rd_data_out[120] rd_data_out[121] rd_data_out[122] rd_data_out[123] rd_data_out[124]
+ rd_data_out[125] rd_data_out[126] rd_data_out[127] rd_data_out[12] rd_data_out[13]
+ rd_data_out[14] rd_data_out[15] rd_data_out[16] rd_data_out[17] rd_data_out[18]
+ rd_data_out[19] rd_data_out[1] rd_data_out[20] rd_data_out[21] rd_data_out[22] rd_data_out[23]
+ rd_data_out[24] rd_data_out[25] rd_data_out[26] rd_data_out[27] rd_data_out[28]
+ rd_data_out[29] rd_data_out[2] rd_data_out[30] rd_data_out[31] rd_data_out[32] rd_data_out[33]
+ rd_data_out[34] rd_data_out[35] rd_data_out[36] rd_data_out[37] rd_data_out[38]
+ rd_data_out[39] rd_data_out[3] rd_data_out[40] rd_data_out[41] rd_data_out[42] rd_data_out[43]
+ rd_data_out[44] rd_data_out[45] rd_data_out[46] rd_data_out[47] rd_data_out[48]
+ rd_data_out[49] rd_data_out[4] rd_data_out[50] rd_data_out[51] rd_data_out[52] rd_data_out[53]
+ rd_data_out[54] rd_data_out[55] rd_data_out[56] rd_data_out[57] rd_data_out[58]
+ rd_data_out[59] rd_data_out[5] rd_data_out[60] rd_data_out[61] rd_data_out[62] rd_data_out[63]
+ rd_data_out[64] rd_data_out[65] rd_data_out[66] rd_data_out[67] rd_data_out[68]
+ rd_data_out[69] rd_data_out[6] rd_data_out[70] rd_data_out[71] rd_data_out[72] rd_data_out[73]
+ rd_data_out[74] rd_data_out[75] rd_data_out[76] rd_data_out[77] rd_data_out[78]
+ rd_data_out[79] rd_data_out[7] rd_data_out[80] rd_data_out[81] rd_data_out[82] rd_data_out[83]
+ rd_data_out[84] rd_data_out[85] rd_data_out[86] rd_data_out[87] rd_data_out[88]
+ rd_data_out[89] rd_data_out[8] rd_data_out[90] rd_data_out[91] rd_data_out[92] rd_data_out[93]
+ rd_data_out[94] rd_data_out[95] rd_data_out[96] rd_data_out[97] rd_data_out[98]
+ rd_data_out[99] rd_data_out[9] read_enable_to_Elpis read_interactive_req_core0 read_value_to_Elpis[0]
+ read_value_to_Elpis[10] read_value_to_Elpis[11] read_value_to_Elpis[12] read_value_to_Elpis[13]
+ read_value_to_Elpis[14] read_value_to_Elpis[15] read_value_to_Elpis[16] read_value_to_Elpis[17]
+ read_value_to_Elpis[18] read_value_to_Elpis[19] read_value_to_Elpis[1] read_value_to_Elpis[20]
+ read_value_to_Elpis[21] read_value_to_Elpis[22] read_value_to_Elpis[23] read_value_to_Elpis[24]
+ read_value_to_Elpis[25] read_value_to_Elpis[26] read_value_to_Elpis[27] read_value_to_Elpis[28]
+ read_value_to_Elpis[29] read_value_to_Elpis[2] read_value_to_Elpis[30] read_value_to_Elpis[31]
+ read_value_to_Elpis[3] read_value_to_Elpis[4] read_value_to_Elpis[5] read_value_to_Elpis[6]
+ read_value_to_Elpis[7] read_value_to_Elpis[8] read_value_to_Elpis[9] ready req_out_core0
+ requested reset_core reset_mem_req rst spare_wen0_to_sram vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] we we_to_sram wr_data[0] wr_data[100] wr_data[101] wr_data[102] wr_data[103]
+ wr_data[104] wr_data[105] wr_data[106] wr_data[107] wr_data[108] wr_data[109] wr_data[10]
+ wr_data[110] wr_data[111] wr_data[112] wr_data[113] wr_data[114] wr_data[115] wr_data[116]
+ wr_data[117] wr_data[118] wr_data[119] wr_data[11] wr_data[120] wr_data[121] wr_data[122]
+ wr_data[123] wr_data[124] wr_data[125] wr_data[126] wr_data[127] wr_data[12] wr_data[13]
+ wr_data[14] wr_data[15] wr_data[16] wr_data[17] wr_data[18] wr_data[19] wr_data[1]
+ wr_data[20] wr_data[21] wr_data[22] wr_data[23] wr_data[24] wr_data[25] wr_data[26]
+ wr_data[27] wr_data[28] wr_data[29] wr_data[2] wr_data[30] wr_data[31] wr_data[32]
+ wr_data[33] wr_data[34] wr_data[35] wr_data[36] wr_data[37] wr_data[38] wr_data[39]
+ wr_data[3] wr_data[40] wr_data[41] wr_data[42] wr_data[43] wr_data[44] wr_data[45]
+ wr_data[46] wr_data[47] wr_data[48] wr_data[49] wr_data[4] wr_data[50] wr_data[51]
+ wr_data[52] wr_data[53] wr_data[54] wr_data[55] wr_data[56] wr_data[57] wr_data[58]
+ wr_data[59] wr_data[5] wr_data[60] wr_data[61] wr_data[62] wr_data[63] wr_data[64]
+ wr_data[65] wr_data[66] wr_data[67] wr_data[68] wr_data[69] wr_data[6] wr_data[70]
+ wr_data[71] wr_data[72] wr_data[73] wr_data[74] wr_data[75] wr_data[76] wr_data[77]
+ wr_data[78] wr_data[79] wr_data[7] wr_data[80] wr_data[81] wr_data[82] wr_data[83]
+ wr_data[84] wr_data[85] wr_data[86] wr_data[87] wr_data[88] wr_data[89] wr_data[8]
+ wr_data[90] wr_data[91] wr_data[92] wr_data[93] wr_data[94] wr_data[95] wr_data[96]
+ wr_data[97] wr_data[98] wr_data[99] wr_data[9]
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2106_ _2149_/CLK _2106_/D vssd1 vssd1 vccd1 vccd1 _2106_/Q sky130_fd_sc_hd__dfxtp_4
X_2037_ _2155_/CLK _2037_/D vssd1 vssd1 vccd1 vccd1 _2037_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1454__A1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1454__B2 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1142__B1 _1958_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1647__754 vssd1 vssd1 vccd1 vccd1 _1647__754/HI la_data_out[95] sky130_fd_sc_hd__conb_1
XANTENNA_input127_A la_data_in[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input92_A la_data_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1381__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output346_A _1686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1270_ _1282_/B vssd1 vssd1 vccd1 vccd1 _1270_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output513_A _2062_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1436__A1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0985_ _0985_/A _0993_/B vssd1 vssd1 vccd1 vccd1 _0986_/A sky130_fd_sc_hd__and2_1
XFILLER_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput401 _1726_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[26] sky130_fd_sc_hd__buf_2
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput434 _1999_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[27] sky130_fd_sc_hd__buf_2
XANTENNA__1057__C _1757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput423 _1959_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[17] sky130_fd_sc_hd__buf_2
Xoutput412 _1707_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[7] sky130_fd_sc_hd__buf_2
Xoutput456 _2126_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[104] sky130_fd_sc_hd__buf_2
Xoutput478 _2146_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[124] sky130_fd_sc_hd__buf_2
XFILLER_114_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput467 _2136_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[114] sky130_fd_sc_hd__buf_2
Xoutput445 _1923_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[8] sky130_fd_sc_hd__buf_2
XFILLER_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1537_ _2101_/Q _1533_/X input59/X _1534_/X vssd1 vssd1 vccd1 vccd1 _2101_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1354__A _2021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput489 _2041_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[19] sky130_fd_sc_hd__buf_2
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1468_ _2021_/Q _1468_/B vssd1 vssd1 vccd1 vccd1 _1507_/A sky130_fd_sc_hd__or2_1
XANTENNA__1073__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1399_ _2134_/Q _1396_/X input60/X _1397_/X vssd1 vssd1 vccd1 vccd1 _2134_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1427__B2 _1425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1427__A1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1963__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1363__B1 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input244_A wr_data[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1418__A1 _2149_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1439__A _1439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2052__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1873__S _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0997__B _1009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output630_A _1122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1322_ _1322_/A _1322_/B vssd1 vssd1 vccd1 vccd1 _1334_/B sky130_fd_sc_hd__or2_1
XFILLER_84_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1253_ _1252_/A _1263_/C _1252_/Y vssd1 vssd1 vccd1 vccd1 _1253_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1184_ _1212_/A _1184_/B vssd1 vssd1 vccd1 vccd1 _1195_/B sky130_fd_sc_hd__or2_1
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1409__A1 _2142_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1349__A _1349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0968_ _0968_/A _0972_/B vssd1 vssd1 vccd1 vccd1 _0969_/A sky130_fd_sc_hd__and2_1
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_133_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1783__S _1922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0899_ _1732_/A _1705_/A vssd1 vssd1 vccd1 vccd1 _0900_/A sky130_fd_sc_hd__and2_1
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1958__S _1958_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2075__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1820__A1 _1688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input194_A wr_data[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input55_A dout0_to_sram[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1722__A _1722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1868__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1940_ _0936_/X _1940_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1940_/X sky130_fd_sc_hd__mux2_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output580_A _1734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1871_ _1870_/X _1331_/Y _2012_/S vssd1 vssd1 vccd1 vccd1 _1871_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1552__659 vssd1 vssd1 vccd1 vccd1 _1552__659/HI la_data_out[0] sky130_fd_sc_hd__conb_1
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1305_ _1305_/A _1305_/B vssd1 vssd1 vccd1 vccd1 _1317_/B sky130_fd_sc_hd__or2_1
XFILLER_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1236_ _1239_/A vssd1 vssd1 vccd1 vccd1 _1244_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1167_ _1168_/B vssd1 vssd1 vccd1 vccd1 _1175_/B sky130_fd_sc_hd__inv_2
XANTENNA__2098__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1098_ _1098_/A vssd1 vssd1 vccd1 vccd1 _1098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1778__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1802__A1 _1685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1079__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_133_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input207_A wr_data[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1717__A _1717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output426_A _1895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2070_ _2155_/CLK _2070_/D vssd1 vssd1 vccd1 vccd1 _2070_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1021_ _1733_/A _2151_/Q _1739_/A vssd1 vssd1 vccd1 vccd1 _1022_/A sky130_fd_sc_hd__and3_1
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ _1922_/X _0912_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1923_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1854_ _1853_/X _1294_/Y _2013_/S vssd1 vssd1 vccd1 vccd1 _1854_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1548__B1 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1785_ _1166_/Y _1784_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1785_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1065__C _1761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1081__B _1081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1219_ _1230_/B vssd1 vssd1 vccd1 vccd1 _1219_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1539__B1 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2113__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1574__681 vssd1 vssd1 vccd1 vccd1 _1574__681/HI la_data_out[22] sky130_fd_sc_hd__conb_1
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1971__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput301 wr_data[92] vssd1 vssd1 vccd1 vccd1 _2000_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input157_A la_data_in[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input18_A addr_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_129_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output543_A _2090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1881__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _2149_/CLK _2122_/D vssd1 vssd1 vccd1 vccd1 _2122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2053_ _2155_/CLK _2053_/D vssd1 vssd1 vccd1 vccd1 _2053_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1004_ _1004_/A vssd1 vssd1 vccd1 vccd1 _1004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2136__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1906_ _1905_/X _1906_/A1 _1938_/S vssd1 vssd1 vccd1 vccd1 _1906_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1558__665 vssd1 vssd1 vccd1 vccd1 _1558__665/HI la_data_out[6] sky130_fd_sc_hd__conb_1
X_1837_ _1836_/X input3/X _1938_/S vssd1 vssd1 vccd1 vccd1 _1837_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1768_ _1142_/Y _1141_/Y _2015_/S vssd1 vssd1 vccd1 vccd1 _1768_/X sky130_fd_sc_hd__mux2_4
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1699_ _1699_/A vssd1 vssd1 vccd1 vccd1 _1699_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1791__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1966__S _2010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_126_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input274_A wr_data[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1267__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput120 la_data_in[52] vssd1 vssd1 vccd1 vccd1 _1720_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput153 la_data_in[82] vssd1 vssd1 vccd1 vccd1 _1752_/A sky130_fd_sc_hd__buf_6
Xinput142 la_data_in[72] vssd1 vssd1 vccd1 vccd1 _1742_/A sky130_fd_sc_hd__buf_6
Xinput131 la_data_in[62] vssd1 vssd1 vccd1 vccd1 _1730_/A sky130_fd_sc_hd__clkbuf_4
Xinput186 wr_data[103] vssd1 vssd1 vccd1 vccd1 _0909_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 la_data_in[92] vssd1 vssd1 vccd1 vccd1 _1762_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput175 read_interactive_req_core0 vssd1 vssd1 vccd1 vccd1 _0857_/A sky130_fd_sc_hd__clkbuf_1
Xinput197 wr_data[113] vssd1 vssd1 vccd1 vccd1 _0951_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1730__A _1730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1999__A0 _1998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output493_A _2044_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1876__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1177__A _1177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput627 _1116_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
Xoutput605 _1737_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[3] sky130_fd_sc_hd__buf_2
Xoutput616 _1096_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput638 _1136_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1484_ _2062_/Q _1479_/X input83/X _1480_/X vssd1 vssd1 vccd1 vccd1 _2062_/D sky130_fd_sc_hd__a22o_1
XFILLER_97_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2105_ _2149_/CLK _2105_/D vssd1 vssd1 vccd1 vccd1 _2105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2036_ _2155_/CLK _2036_/D vssd1 vssd1 vccd1 vccd1 _2036_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1454__A2 _1452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1786__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1087__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input85_A la_data_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1725__A _1725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1381__A1 _2122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output339_A _1698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output506_A _2056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_repeater656_A _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0984_ _0984_/A vssd1 vssd1 vccd1 vccd1 _0984_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput402 _1727_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[27] sky130_fd_sc_hd__buf_2
Xoutput424 _1963_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[18] sky130_fd_sc_hd__buf_2
XFILLER_114_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput435 _2003_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[28] sky130_fd_sc_hd__buf_2
Xoutput413 _1708_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[8] sky130_fd_sc_hd__buf_2
Xoutput468 _2137_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[115] sky130_fd_sc_hd__buf_2
X_1536_ _2100_/Q _1533_/X input58/X _1534_/X vssd1 vssd1 vccd1 vccd1 _2100_/D sky130_fd_sc_hd__a22o_1
Xoutput457 _2127_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[105] sky130_fd_sc_hd__buf_2
Xoutput446 _1927_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[9] sky130_fd_sc_hd__buf_2
Xoutput479 _2147_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[125] sky130_fd_sc_hd__buf_2
XFILLER_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1467_ input77/X _1438_/A _2053_/Q _1439_/A vssd1 vssd1 vccd1 vccd1 _2053_/D sky130_fd_sc_hd__o22a_1
XANTENNA__1073__C _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1398_ _2133_/Q _1396_/X input59/X _1397_/X vssd1 vssd1 vccd1 vccd1 _2133_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1370__A _2020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2019_ _2155_/CLK _2019_/D vssd1 vssd1 vccd1 vccd1 _2019_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__1427__A2 _1422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1614__721 vssd1 vssd1 vccd1 vccd1 _1614__721/HI la_data_out[62] sky130_fd_sc_hd__conb_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1363__A1 _2113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input237_A wr_data[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1280__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output456_A _2126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output623_A _1110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1321_ _1319_/C _1308_/X _1320_/Y vssd1 vssd1 vccd1 vccd1 _1321_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1252_ _1252_/A _1263_/C vssd1 vssd1 vccd1 vccd1 _1252_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1183_ _1212_/A _1182_/B _1193_/B vssd1 vssd1 vccd1 vccd1 _1183_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0967_ _0967_/A vssd1 vssd1 vccd1 vccd1 _0967_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0898_ _0898_/A vssd1 vssd1 vccd1 vccd1 _0898_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1519_ _1519_/A vssd1 vssd1 vccd1 vccd1 _1519_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1974__S _1990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input187_A wr_data[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input48_A core0_data_print[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1870_ input9/X _1333_/X _1882_/S vssd1 vssd1 vccd1 vccd1 _1870_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output573_A _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1884__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1591__698 vssd1 vssd1 vccd1 vccd1 _1591__698/HI la_data_out[39] sky130_fd_sc_hd__conb_1
XFILLER_123_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1304_ input7/X _1293_/Y _1314_/B vssd1 vssd1 vccd1 vccd1 _1304_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1235_ _1235_/A vssd1 vssd1 vccd1 vccd1 _1239_/A sky130_fd_sc_hd__inv_2
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1166_ _1175_/A _1175_/C _1165_/Y vssd1 vssd1 vccd1 vccd1 _1166_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1097_ _2019_/Q _1097_/B vssd1 vssd1 vccd1 vccd1 _1098_/A sky130_fd_sc_hd__and2_1
XFILLER_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1794__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1999_ _1998_/X _0992_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1999_/X sky130_fd_sc_hd__mux2_4
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1095__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1318__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2042__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1969__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input102_A la_data_in[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0902__A _0902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_125_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1309__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1733__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output321_A _1779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1020_ _1020_/A vssd1 vssd1 vccd1 vccd1 _1020_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1879__S _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1922_ _1921_/X _1922_/A1 _1922_/S vssd1 vssd1 vccd1 vccd1 _1922_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1796__A1 _1684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1853_ _1852_/X _1296_/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1853_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1548__A1 _2110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1784_ _1783_/X _1682_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1784_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2065__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1218_ _1218_/A _1218_/B vssd1 vssd1 vccd1 vccd1 _1230_/B sky130_fd_sc_hd__or2_1
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1789__S _1922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1484__B1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1149_ _0875_/A _1144_/X _1148_/Y vssd1 vssd1 vccd1 vccd1 _1149_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1539__B2 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput302 wr_data[93] vssd1 vssd1 vccd1 vccd1 _2004_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1475__B1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1728__A _1728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_113_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2088__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1950__A1 _1950_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output536_A _2083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2121_ _2149_/CLK _2121_/D vssd1 vssd1 vccd1 vccd1 _2121_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2052_ _2155_/CLK _2052_/D vssd1 vssd1 vccd1 vccd1 _2052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1003_ _1732_/A _1730_/A vssd1 vssd1 vccd1 vccd1 _1004_/A sky130_fd_sc_hd__and2_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1905_ _1904_/X _1905_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1905_/X sky130_fd_sc_hd__mux2_4
X_1836_ _1835_/X _1259_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1836_/X sky130_fd_sc_hd__mux2_1
X_1767_ _1767_/A0 _1767_/A1 _1767_/S vssd1 vssd1 vccd1 vccd1 _1767_/X sky130_fd_sc_hd__mux2_8
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1698_ _1698_/A vssd1 vssd1 vccd1 vccd1 _1698_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_106_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1457__B1 _2045_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1982__S _2010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input267_A wr_data[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput110 la_data_in[43] vssd1 vssd1 vccd1 vccd1 _1711_/A sky130_fd_sc_hd__buf_4
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput121 la_data_in[53] vssd1 vssd1 vccd1 vccd1 _1721_/A sky130_fd_sc_hd__buf_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input30_A core0_data_print[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput132 la_data_in[63] vssd1 vssd1 vccd1 vccd1 _1731_/A sky130_fd_sc_hd__buf_6
Xinput143 la_data_in[73] vssd1 vssd1 vccd1 vccd1 _1743_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput154 la_data_in[83] vssd1 vssd1 vccd1 vccd1 _1753_/A sky130_fd_sc_hd__clkbuf_2
Xinput165 la_data_in[93] vssd1 vssd1 vccd1 vccd1 _1763_/A sky130_fd_sc_hd__buf_2
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput187 wr_data[104] vssd1 vssd1 vccd1 vccd1 _0914_/A sky130_fd_sc_hd__buf_2
Xinput176 req_out_core0 vssd1 vssd1 vccd1 vccd1 _0861_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput198 wr_data[114] vssd1 vssd1 vccd1 vccd1 _0956_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1448__B1 _2038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output486_A _2038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput617 _1098_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XANTENNA__1892__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput606 _1738_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[4] sky130_fd_sc_hd__buf_2
Xoutput639 _1138_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_99_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput628 _1118_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
X_1631__738 vssd1 vssd1 vccd1 vccd1 _1631__738/HI la_data_out[79] sky130_fd_sc_hd__conb_1
X_1483_ _2061_/Q _1479_/X input82/X _1480_/X vssd1 vssd1 vccd1 vccd1 _2061_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2104_ _2149_/CLK _2104_/D vssd1 vssd1 vccd1 vccd1 _2104_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2103__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2035_ _2155_/CLK _2035_/D vssd1 vssd1 vccd1 vccd1 _2035_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1819_ _1818_/X _1223_/A _1938_/S vssd1 vssd1 vccd1 vccd1 _1819_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1914__A1 _1914_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1977__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_127_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input78_A dout0_to_sram[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1905__A1 _1905_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2126__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1741__A _1741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1887__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater649_A _1942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0983_ _1732_/A _1725_/A vssd1 vssd1 vccd1 vccd1 _0984_/A sky130_fd_sc_hd__and2_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput425 _1967_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[19] sky130_fd_sc_hd__buf_2
Xoutput403 _1728_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[28] sky130_fd_sc_hd__buf_2
Xoutput414 _1709_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[9] sky130_fd_sc_hd__buf_2
Xoutput436 _2007_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[29] sky130_fd_sc_hd__buf_2
Xoutput458 _2128_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[106] sky130_fd_sc_hd__buf_2
XFILLER_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1535_ _2099_/Q _1533_/X input57/X _1534_/X vssd1 vssd1 vccd1 vccd1 _2099_/D sky130_fd_sc_hd__a22o_1
Xoutput447 _1732_/X vssd1 vssd1 vccd1 vccd1 is_loading_memory_into_core sky130_fd_sc_hd__buf_2
Xoutput469 _2138_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[116] sky130_fd_sc_hd__buf_2
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1466_ input76/X _1438_/A _2052_/Q _1439_/A vssd1 vssd1 vccd1 vccd1 _2052_/D sky130_fd_sc_hd__o22a_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1397_ _1411_/A vssd1 vssd1 vccd1 vccd1 _1397_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ _2155_/CLK _2018_/D vssd1 vssd1 vccd1 vccd1 _2018_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1797__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1653__760 vssd1 vssd1 vccd1 vccd1 _1653__760/HI la_data_out[102] sky130_fd_sc_hd__conb_1
XANTENNA__2149__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input132_A la_data_in[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0905__A _0905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1736__A _1736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output351_A _1012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1320_ _1343_/C vssd1 vssd1 vccd1 vccd1 _1320_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1251_ input2/X _1240_/Y _1260_/B vssd1 vssd1 vccd1 vccd1 _1251_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1182_ _1186_/A _1182_/B vssd1 vssd1 vccd1 vccd1 _1193_/B sky130_fd_sc_hd__or2_1
XFILLER_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1596__703 vssd1 vssd1 vccd1 vccd1 _1596__703/HI la_data_out[44] sky130_fd_sc_hd__conb_1
XANTENNA__1290__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0966_ _1732_/A _1721_/A vssd1 vssd1 vccd1 vccd1 _0967_/A sky130_fd_sc_hd__and2_1
X_1637__744 vssd1 vssd1 vccd1 vccd1 _1637__744/HI la_data_out[85] sky130_fd_sc_hd__conb_1
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0897_ _0897_/A _0909_/B vssd1 vssd1 vccd1 vccd1 _0898_/A sky130_fd_sc_hd__and2_2
XFILLER_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1518_ _2088_/Q _1366_/X input75/X _1367_/X vssd1 vssd1 vccd1 vccd1 _2088_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1449_ input61/X _1445_/X _2039_/Q _1446_/X vssd1 vssd1 vccd1 vccd1 _2039_/D sky130_fd_sc_hd__o22a_1
XFILLER_56_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1990__S _1990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1291__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output399_A _1724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output566_A _2111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1303_ _1303_/A _1319_/B vssd1 vssd1 vccd1 vccd1 _1314_/B sky130_fd_sc_hd__or2_1
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1234_ _1232_/A _1232_/B _1233_/Y vssd1 vssd1 vccd1 vccd1 _1234_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1165_ _1175_/A _1175_/C vssd1 vssd1 vccd1 vccd1 _1165_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1096_ _1096_/A vssd1 vssd1 vccd1 vccd1 _1096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1998_ _1997_/X _1998_/A1 _2014_/S vssd1 vssd1 vccd1 vccd1 _1998_/X sky130_fd_sc_hd__mux2_2
XFILLER_119_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0949_ _1732_/A _1717_/A vssd1 vssd1 vccd1 vccd1 _0950_/A sky130_fd_sc_hd__and2_1
XFILLER_134_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1985__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input297_A wr_data[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input60_A dout0_to_sram[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1921_ _1920_/X _1921_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1921_/X sky130_fd_sc_hd__mux2_2
XANTENNA__1895__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1245__A1 _1235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1852_ input6/X _1298_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1852_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1783_ _1782_/X _1168_/A _1922_/S vssd1 vssd1 vccd1 vccd1 _1783_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1217_ _1218_/A _1215_/B _1216_/Y vssd1 vssd1 vccd1 vccd1 _1217_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1484__A1 _2062_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1148_ _1148_/A _1152_/A vssd1 vssd1 vccd1 vccd1 _1148_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1079_ _2019_/Q _1079_/B vssd1 vssd1 vccd1 vccd1 _1080_/A sky130_fd_sc_hd__and2_1
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1539__A2 _1533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput303 wr_data[94] vssd1 vssd1 vccd1 vccd1 _2008_/A1 sky130_fd_sc_hd__buf_2
XFILLER_102_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1475__A1 _2055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input212_A wr_data[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1475__B2 _1473_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1744__A _1744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output529_A _2077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output431_A _1987_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2120_ _2149_/CLK _2120_/D vssd1 vssd1 vccd1 vccd1 _2120_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2051_ _2155_/CLK _2051_/D vssd1 vssd1 vccd1 vccd1 _2051_/Q sky130_fd_sc_hd__dfxtp_2
X_1002_ _1002_/A vssd1 vssd1 vccd1 vccd1 _1002_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1466__B2 _1439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1466__A1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1904_ _0898_/X _1904_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1904_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1835_ _1834_/X _1262_/Y _2012_/S vssd1 vssd1 vccd1 vccd1 _1835_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2032__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1766_ _1766_/A vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1697_ _1697_/A vssd1 vssd1 vccd1 vccd1 _1697_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1457__A1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1457__B2 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1393__B1 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input162_A la_data_in[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput111 la_data_in[44] vssd1 vssd1 vccd1 vccd1 _1712_/A sky130_fd_sc_hd__buf_6
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput100 la_data_in[34] vssd1 vssd1 vccd1 vccd1 _1702_/A sky130_fd_sc_hd__buf_2
XFILLER_103_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput144 la_data_in[74] vssd1 vssd1 vccd1 vccd1 _1744_/A sky130_fd_sc_hd__buf_2
Xinput133 la_data_in[64] vssd1 vssd1 vccd1 vccd1 _1734_/A sky130_fd_sc_hd__clkbuf_1
Xinput122 la_data_in[54] vssd1 vssd1 vccd1 vccd1 _1722_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput155 la_data_in[84] vssd1 vssd1 vccd1 vccd1 _1754_/A sky130_fd_sc_hd__buf_6
XANTENNA_input23_A core0_data_print[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput166 la_data_in[94] vssd1 vssd1 vccd1 vccd1 _1764_/A sky130_fd_sc_hd__buf_6
XFILLER_102_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput177 requested vssd1 vssd1 vccd1 vccd1 _0866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput188 wr_data[105] vssd1 vssd1 vccd1 vccd1 _0918_/A sky130_fd_sc_hd__clkbuf_1
Xinput199 wr_data[115] vssd1 vssd1 vccd1 vccd1 _0960_/A sky130_fd_sc_hd__buf_4
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1448__A1 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1739__A _1739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2055__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output381_A _1028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output479_A _2147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput607 _1739_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[5] sky130_fd_sc_hd__buf_2
Xoutput618 _1100_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XANTENNA__1384__B1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput629 _1120_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
X_1670__777 vssd1 vssd1 vccd1 vccd1 _1670__777/HI la_data_out[119] sky130_fd_sc_hd__conb_1
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1482_ _2060_/Q _1479_/X input81/X _1480_/X vssd1 vssd1 vccd1 vccd1 _2060_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2103_ _1767_/X _2103_/D vssd1 vssd1 vccd1 vccd1 _2103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2034_ _2155_/CLK _2034_/D vssd1 vssd1 vccd1 vccd1 _2034_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1564__671 vssd1 vssd1 vccd1 vccd1 _1564__671/HI la_data_out[12] sky130_fd_sc_hd__conb_1
XFILLER_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1818_ _1817_/X _1227_/Y _2013_/S vssd1 vssd1 vccd1 vccd1 _1818_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_117_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_116_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1749_ _1749_/A vssd1 vssd1 vccd1 vccd1 _1749_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2078__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1850__A1 _1693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1993__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0982_ _0982_/A vssd1 vssd1 vccd1 vccd1 _0982_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput426 _1895_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[1] sky130_fd_sc_hd__buf_2
Xoutput415 _1891_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[0] sky130_fd_sc_hd__buf_2
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput404 _1729_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[29] sky130_fd_sc_hd__buf_2
Xoutput459 _2129_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[107] sky130_fd_sc_hd__buf_2
Xoutput437 _1899_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[2] sky130_fd_sc_hd__buf_2
XFILLER_114_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1534_ _1541_/A vssd1 vssd1 vccd1 vccd1 _1534_/X sky130_fd_sc_hd__buf_2
XFILLER_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput448 _0859_/X vssd1 vssd1 vccd1 vccd1 is_ready_dataout_core0 sky130_fd_sc_hd__buf_2
XFILLER_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1465_ input74/X _1459_/X _2051_/Q _1460_/X vssd1 vssd1 vccd1 vccd1 _2051_/D sky130_fd_sc_hd__o22a_1
X_1396_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1396_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2017_ _0875_/A _0866_/A _2017_/S vssd1 vssd1 vccd1 vccd1 _2017_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input125_A la_data_in[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1988__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0905__B _0909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input90_A la_data_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_127_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2000__A1 _2000_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1752__A _1752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1250_ _1263_/A _1250_/B vssd1 vssd1 vccd1 vccd1 _1260_/B sky130_fd_sc_hd__or2_1
XFILLER_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output511_A _2061_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1181_ _1177_/A _1179_/A _1191_/B vssd1 vssd1 vccd1 vccd1 _1181_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1511__B1 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output609_A _1741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1898__S _1934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1814__A1 _1687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_119_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0965_ _0965_/A vssd1 vssd1 vccd1 vccd1 _0965_/X sky130_fd_sc_hd__clkbuf_1
X_1676__783 vssd1 vssd1 vccd1 vccd1 _1676__783/HI la_data_out[125] sky130_fd_sc_hd__conb_1
X_0896_ _0896_/A vssd1 vssd1 vccd1 vccd1 _0896_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1517_ _2087_/Q _1366_/X input64/X _1367_/X vssd1 vssd1 vccd1 vccd1 _2087_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1448_ input60/X _1445_/X _2038_/Q _1446_/X vssd1 vssd1 vccd1 vccd1 _2038_/D sky130_fd_sc_hd__o22a_1
XFILLER_4_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1379_ _2120_/Q _1373_/X input75/X _1376_/X vssd1 vssd1 vccd1 vccd1 _2120_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1502__B1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__2116__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input242_A wr_data[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0916__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1747__A _1747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output461_A _2131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output559_A _2104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1302_ _1302_/A _1305_/A vssd1 vssd1 vccd1 vccd1 _1319_/B sky130_fd_sc_hd__or2_1
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1233_ _1244_/B vssd1 vssd1 vccd1 vccd1 _1233_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1164_ _2152_/Q _1150_/A _1148_/Y _1155_/X vssd1 vssd1 vccd1 vccd1 _1175_/C sky130_fd_sc_hd__a22oi_2
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1095_ _2019_/Q _1095_/B vssd1 vssd1 vccd1 vccd1 _1096_/A sky130_fd_sc_hd__and2_1
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1604__711 vssd1 vssd1 vccd1 vccd1 _1604__711/HI la_data_out[52] sky130_fd_sc_hd__conb_1
XANTENNA__2139__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ _1996_/X _1997_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1997_/X sky130_fd_sc_hd__mux2_1
X_0948_ _0948_/A vssd1 vssd1 vccd1 vccd1 _0948_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0879_ _0879_/A _1882_/S vssd1 vssd1 vccd1 vccd1 _0880_/A sky130_fd_sc_hd__and2_1
XANTENNA__1971__A0 _1970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input192_A wr_data[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input53_A dout0_to_sram[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1920_ _0915_/X _1920_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1920_/X sky130_fd_sc_hd__mux2_4
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1851_ _1290_/X _1850_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1851_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1782_ _1781_/X _1158_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1782_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1953__A0 _1952_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1181__A1 _1177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1216_ _1228_/B vssd1 vssd1 vccd1 vccd1 _1216_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1147_ _1147_/A vssd1 vssd1 vccd1 vccd1 _1887_/S sky130_fd_sc_hd__buf_12
XFILLER_26_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1078_ _1078_/A vssd1 vssd1 vccd1 vccd1 _1078_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_107_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_134_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput304 wr_data[95] vssd1 vssd1 vccd1 vccd1 _2012_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1475__A2 _1470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1996__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input205_A wr_data[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1581__688 vssd1 vssd1 vccd1 vccd1 _1581__688/HI la_data_out[29] sky130_fd_sc_hd__conb_1
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output424_A _1963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1760__A _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2050_ _2155_/CLK _2050_/D vssd1 vssd1 vccd1 vccd1 _2050_/Q sky130_fd_sc_hd__dfxtp_2
X_1001_ _1001_/A _1009_/B vssd1 vssd1 vccd1 vccd1 _1002_/A sky130_fd_sc_hd__and2_1
XFILLER_75_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1466__A2 _1438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1903_ _1902_/X _0890_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1903_/X sky130_fd_sc_hd__mux2_2
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1834_ input3/X _1264_/X _1882_/S vssd1 vssd1 vccd1 vccd1 _1834_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1765_ _1765_/A vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__buf_2
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1696_ _1696_/A vssd1 vssd1 vccd1 vccd1 _1696_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1457__A2 _1452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1917__A0 _1916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1393__A1 _2130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input155_A la_data_in[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput101 la_data_in[35] vssd1 vssd1 vccd1 vccd1 _1703_/A sky130_fd_sc_hd__buf_4
XFILLER_49_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput145 la_data_in[75] vssd1 vssd1 vccd1 vccd1 _1745_/A sky130_fd_sc_hd__buf_8
XFILLER_103_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput134 la_data_in[65] vssd1 vssd1 vccd1 vccd1 _1735_/A sky130_fd_sc_hd__buf_4
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput112 la_data_in[45] vssd1 vssd1 vccd1 vccd1 _1713_/A sky130_fd_sc_hd__buf_4
Xinput123 la_data_in[55] vssd1 vssd1 vccd1 vccd1 _1723_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1145__B2 _0876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput156 la_data_in[85] vssd1 vssd1 vccd1 vccd1 _1755_/A sky130_fd_sc_hd__clkbuf_2
Xinput167 la_data_in[95] vssd1 vssd1 vccd1 vccd1 _1765_/A sky130_fd_sc_hd__buf_4
Xinput178 reset_mem_req vssd1 vssd1 vccd1 vccd1 _0843_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA_input16_A addr_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput189 wr_data[106] vssd1 vssd1 vccd1 vccd1 _0922_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_112_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0924__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput608 _1740_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[6] sky130_fd_sc_hd__buf_2
XFILLER_126_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1755__A _1755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1550_ _0870_/A _0841_/X _2155_/Q _1549_/Y _0852_/B vssd1 vssd1 vccd1 vccd1 _2155_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__1384__A1 _2123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput619 _1102_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA_output639_A _1138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output541_A _2088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1481_ _2059_/Q _1479_/X input80/X _1480_/X vssd1 vssd1 vccd1 vccd1 _2059_/D sky130_fd_sc_hd__a22o_1
XFILLER_121_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2102_ _2149_/CLK _2102_/D vssd1 vssd1 vccd1 vccd1 _2102_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2033_ _2155_/CLK _2033_/D vssd1 vssd1 vccd1 vccd1 _2033_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1817_ _1816_/X _1229_/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1817_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1748_ _1748_/A vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A addr_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input272_A wr_data[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0919__A _0919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1587__694 vssd1 vssd1 vccd1 vccd1 _1587__694/HI la_data_out[35] sky130_fd_sc_hd__conb_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2022__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output491_A _2042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0981_ _0981_/A _0993_/B vssd1 vssd1 vccd1 vccd1 _0982_/A sky130_fd_sc_hd__and2_1
XFILLER_60_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput405 _1702_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[2] sky130_fd_sc_hd__buf_2
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput416 _1931_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[10] sky130_fd_sc_hd__buf_2
XFILLER_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1533_ _1540_/A vssd1 vssd1 vccd1 vccd1 _1533_/X sky130_fd_sc_hd__buf_2
Xoutput438 _2011_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[30] sky130_fd_sc_hd__buf_2
Xoutput427 _1971_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[20] sky130_fd_sc_hd__buf_2
Xoutput449 _1419_/A vssd1 vssd1 vccd1 vccd1 is_ready_print_core0 sky130_fd_sc_hd__buf_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1464_ input73/X _1459_/X _2050_/Q _1460_/X vssd1 vssd1 vccd1 vccd1 _2050_/D sky130_fd_sc_hd__o22a_1
XFILLER_86_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1395_ _2132_/Q _1389_/X input58/X _1390_/X vssd1 vssd1 vccd1 vccd1 _2132_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2016_ _1766_/A _2016_/A1 _2016_/S vssd1 vssd1 vccd1 vccd1 _2016_/X sky130_fd_sc_hd__mux2_2
XFILLER_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_128_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2045__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A la_data_in[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1621__728 vssd1 vssd1 vccd1 vccd1 _1621__728/HI la_data_out[69] sky130_fd_sc_hd__conb_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input83_A dout0_to_sram[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output337_A _1696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1180_ _1212_/A _1213_/D vssd1 vssd1 vccd1 vccd1 _1191_/B sky130_fd_sc_hd__or2_1
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1511__A1 _2081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater654_A _1958_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0964_ _0964_/A _0972_/B vssd1 vssd1 vccd1 vccd1 _0965_/A sky130_fd_sc_hd__and2_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0895_ _1732_/A _1704_/A vssd1 vssd1 vccd1 vccd1 _0896_/A sky130_fd_sc_hd__and2_1
XFILLER_134_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1516_ _2086_/Q _1366_/X input53/X _1367_/X vssd1 vssd1 vccd1 vccd1 _2086_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2068__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1447_ input59/X _1445_/X _2037_/Q _1446_/X vssd1 vssd1 vccd1 vccd1 _2037_/D sky130_fd_sc_hd__o22a_1
X_1378_ _2119_/Q _1373_/X input64/X _1376_/X vssd1 vssd1 vccd1 vccd1 _2119_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1502__A1 _2074_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input235_A wr_data[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1999__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0932__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_127_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1980__A1 _1980_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1763__A _1763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output454_A _2124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output621_A _1106_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1301_ input7/X vssd1 vssd1 vccd1 vccd1 _1305_/A sky130_fd_sc_hd__inv_2
X_1232_ _1232_/A _1232_/B vssd1 vssd1 vccd1 vccd1 _1244_/B sky130_fd_sc_hd__or2_1
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1496__B1 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1163_ _1144_/X _1160_/A _1175_/A _1162_/X vssd1 vssd1 vccd1 vccd1 _1163_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1094_ _1094_/A vssd1 vssd1 vccd1 vccd1 _1094_/X sky130_fd_sc_hd__clkbuf_1
X_1643__750 vssd1 vssd1 vccd1 vccd1 _1643__750/HI la_data_out[91] sky130_fd_sc_hd__conb_1
XFILLER_100_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1003__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1996_ _0994_/X _1996_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1996_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0947_ _0947_/A _0951_/B vssd1 vssd1 vccd1 vccd1 _0948_/A sky130_fd_sc_hd__and2_1
XFILLER_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0878_ _0976_/A vssd1 vssd1 vccd1 vccd1 _1882_/S sky130_fd_sc_hd__buf_12
XFILLER_106_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_71_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_137_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_137_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input185_A wr_data[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1962__A1 _1962_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input46_A core0_data_print[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1478__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1627__734 vssd1 vssd1 vccd1 vccd1 _1627__734/HI la_data_out[75] sky130_fd_sc_hd__conb_1
XFILLER_34_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1758__A _1758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1850_ _1849_/X _1693_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1850_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output571_A _2115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1781_ _1780_/X _1161_/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1781_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1402__B1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1953__A1 _1953_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_112_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2106__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1215_ _1218_/A _1215_/B vssd1 vssd1 vccd1 vccd1 _1228_/B sky130_fd_sc_hd__or2_1
XFILLER_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1146_ _1732_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _1147_/A sky130_fd_sc_hd__or2_1
XFILLER_1_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1077_ _2019_/Q _1077_/B vssd1 vssd1 vccd1 vccd1 _1078_/A sky130_fd_sc_hd__and2_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1979_ _1978_/X _0971_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1979_/X sky130_fd_sc_hd__mux2_2
XFILLER_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_134_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput305 wr_data[96] vssd1 vssd1 vccd1 vccd1 _0879_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1172__A2 _1150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input100_A la_data_in[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2129__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output417_A _1935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1000_ _1000_/A vssd1 vssd1 vccd1 vccd1 _1000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ _1901_/X _1902_/A1 _1958_/S vssd1 vssd1 vccd1 vccd1 _1902_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1833_ _1256_/Y _1832_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1833_/X sky130_fd_sc_hd__mux2_4
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1764_ _1764_/A vssd1 vssd1 vccd1 vccd1 _1764_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1926__A1 _1926_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1695_ _1695_/A vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1129_ _2019_/Q _1129_/B vssd1 vssd1 vccd1 vccd1 _1130_/A sky130_fd_sc_hd__and2_1
XFILLER_14_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1917__A1 _1917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput102 la_data_in[36] vssd1 vssd1 vccd1 vccd1 _1704_/A sky130_fd_sc_hd__buf_6
XANTENNA__1145__A2 _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input148_A la_data_in[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput135 la_data_in[66] vssd1 vssd1 vccd1 vccd1 _1736_/A sky130_fd_sc_hd__buf_8
XFILLER_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput113 la_data_in[46] vssd1 vssd1 vccd1 vccd1 _1714_/A sky130_fd_sc_hd__buf_2
Xinput124 la_data_in[56] vssd1 vssd1 vccd1 vccd1 _1724_/A sky130_fd_sc_hd__buf_2
Xinput146 la_data_in[76] vssd1 vssd1 vccd1 vccd1 _1746_/A sky130_fd_sc_hd__clkbuf_4
Xinput168 la_data_in[96] vssd1 vssd1 vccd1 vccd1 _1767_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput157 la_data_in[86] vssd1 vssd1 vccd1 vccd1 _1756_/A sky130_fd_sc_hd__buf_4
XFILLER_57_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput179 wb_clk_i vssd1 vssd1 vccd1 vccd1 _1767_/A1 sky130_fd_sc_hd__buf_8
XFILLER_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1800__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0924__B _1711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1101__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_126_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1908__A1 _1908_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput609 _1741_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[7] sky130_fd_sc_hd__buf_2
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1480_ _1487_/A vssd1 vssd1 vccd1 vccd1 _1480_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output534_A _2027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2101_ _2149_/CLK _2101_/D vssd1 vssd1 vccd1 vccd1 _2101_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2032_ _2155_/CLK _2032_/D vssd1 vssd1 vccd1 vccd1 _2032_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1011__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1816_ _1223_/A _1231_/X _1882_/S vssd1 vssd1 vccd1 vccd1 _1816_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1747_ _1747_/A vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input265_A wr_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0935__A _0935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0980_ _0980_/A vssd1 vssd1 vccd1 vccd1 _0980_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output484_A _2036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1766__A _1766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput417 _1935_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[11] sky130_fd_sc_hd__buf_2
Xoutput406 _1730_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[30] sky130_fd_sc_hd__buf_2
Xoutput439 _2015_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[31] sky130_fd_sc_hd__buf_2
XFILLER_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1532_ _2098_/Q _1526_/X input56/X _1527_/X vssd1 vssd1 vccd1 vccd1 _2098_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput428 _1975_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[21] sky130_fd_sc_hd__buf_2
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1463_ input72/X _1459_/X _2049_/Q _1460_/X vssd1 vssd1 vccd1 vccd1 _2049_/D sky130_fd_sc_hd__o22a_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1394_ _2131_/Q _1389_/X input57/X _1390_/X vssd1 vssd1 vccd1 vccd1 _2131_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1006__A _1006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2015_ _2014_/X _1008_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _2015_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1660__767 vssd1 vssd1 vccd1 vccd1 _1660__767/HI la_data_out[109] sky130_fd_sc_hd__conb_1
XFILLER_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input76_A dout0_to_sram[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1554__661 vssd1 vssd1 vccd1 vccd1 _1554__661/HI la_data_out[2] sky130_fd_sc_hd__conb_1
XFILLER_135_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0963_ _0963_/A vssd1 vssd1 vccd1 vccd1 _0963_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0894_ _0894_/A vssd1 vssd1 vccd1 vccd1 _0894_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1515_ _2085_/Q _1486_/A input77/X _1487_/A vssd1 vssd1 vccd1 vccd1 _2085_/D sky130_fd_sc_hd__a22o_1
XFILLER_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1446_ _1460_/A vssd1 vssd1 vccd1 vccd1 _1446_/X sky130_fd_sc_hd__clkbuf_2
X_1377_ _2118_/Q _1373_/X input53/X _1376_/X vssd1 vssd1 vccd1 vccd1 _2118_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1266__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input130_A la_data_in[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input228_A wr_data[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0932__B _1713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1300_ _1297_/A _1310_/A _1299_/Y vssd1 vssd1 vccd1 vccd1 _1300_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1231_ _1223_/A _1219_/Y _1242_/B vssd1 vssd1 vccd1 vccd1 _1231_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1496__A1 _2070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1162_ input1/X _1150_/A _1168_/A vssd1 vssd1 vccd1 vccd1 _1162_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1093_ _2019_/Q _1093_/B vssd1 vssd1 vccd1 vccd1 _1094_/A sky130_fd_sc_hd__and2_1
XFILLER_64_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1003__B _1730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1995_ _1994_/X _0988_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1995_/X sky130_fd_sc_hd__mux2_4
XFILLER_119_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2035__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0946_ _0946_/A vssd1 vssd1 vccd1 vccd1 _0946_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0877_ _0891_/A vssd1 vssd1 vccd1 vccd1 _0976_/A sky130_fd_sc_hd__buf_2
XFILLER_133_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1429_ input78/X _1422_/X _2025_/Q _1425_/X vssd1 vssd1 vccd1 vccd1 _2025_/D sky130_fd_sc_hd__o22a_1
XFILLER_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_34_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_7_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_137_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_137_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input178_A reset_mem_req vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input39_A core0_data_print[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1803__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1666__773 vssd1 vssd1 vccd1 vccd1 _1666__773/HI la_data_out[115] sky130_fd_sc_hd__conb_1
XANTENNA__1478__B2 _1473_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0943__A _0943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2058__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output397_A _1722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1780_ _1168_/A _1163_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1780_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1402__A1 _2137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output564_A _2109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1402__B2 _1397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1214_ _1210_/A _1202_/Y _1225_/B vssd1 vssd1 vccd1 vccd1 _1214_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1145_ input1/X _1882_/S _1144_/X _0876_/A vssd1 vssd1 vccd1 vccd1 _1145_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1076_ _1076_/A vssd1 vssd1 vccd1 vccd1 _1076_/X sky130_fd_sc_hd__buf_4
XFILLER_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1978_ _1977_/X _1978_/A1 _2014_/S vssd1 vssd1 vccd1 vccd1 _1978_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1684__A _1684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0929_ _0929_/A vssd1 vssd1 vccd1 vccd1 _0929_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput306 wr_data[97] vssd1 vssd1 vccd1 vccd1 _0883_/A sky130_fd_sc_hd__buf_2
XFILLER_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1880__A1 _1698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input295_A wr_data[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output312_A _1839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1901_ _1900_/X _1901_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1901_/X sky130_fd_sc_hd__mux2_8
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1832_ _1831_/X _1690_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1832_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1763_ _1763_/A vssd1 vssd1 vccd1 vccd1 _1763_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1387__B1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1694_ _1694_/A vssd1 vssd1 vccd1 vccd1 _1694_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1009__A _1009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1128_ _1128_/A vssd1 vssd1 vccd1 vccd1 _1128_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1862__A1 _1695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1059_ _1733_/A _2151_/Q _1758_/A vssd1 vssd1 vccd1 vccd1 _1060_/A sky130_fd_sc_hd__and3_1
XFILLER_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1378__B1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput114 la_data_in[47] vssd1 vssd1 vccd1 vccd1 _1715_/A sky130_fd_sc_hd__buf_2
Xinput103 la_data_in[37] vssd1 vssd1 vccd1 vccd1 _1705_/A sky130_fd_sc_hd__buf_6
XFILLER_103_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput136 la_data_in[67] vssd1 vssd1 vccd1 vccd1 _1737_/A sky130_fd_sc_hd__clkbuf_4
Xinput125 la_data_in[57] vssd1 vssd1 vccd1 vccd1 _1725_/A sky130_fd_sc_hd__buf_4
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput147 la_data_in[77] vssd1 vssd1 vccd1 vccd1 _1747_/A sky130_fd_sc_hd__buf_4
XFILLER_102_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput158 la_data_in[87] vssd1 vssd1 vccd1 vccd1 _1757_/A sky130_fd_sc_hd__clkbuf_2
Xinput169 la_data_in[97] vssd1 vssd1 vccd1 vccd1 _1766_/A sky130_fd_sc_hd__buf_4
XFILLER_91_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input210_A wr_data[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input308_A wr_data[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1101__B _1101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1369__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output527_A _2075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2100_ _2149_/CLK _2100_/D vssd1 vssd1 vccd1 vccd1 _2100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2031_ _2155_/CLK _2031_/D vssd1 vssd1 vccd1 vccd1 _2031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1844__A1 _1692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1011__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1815_ _1222_/X _1814_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1815_/X sky130_fd_sc_hd__mux2_8
X_1746_ _1746_/A vssd1 vssd1 vccd1 vccd1 _1746_/X sky130_fd_sc_hd__buf_4
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1571__678 vssd1 vssd1 vccd1 vccd1 _1571__678/HI la_data_out[19] sky130_fd_sc_hd__conb_1
XFILLER_131_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1532__B1 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1901__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2119__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input160_A la_data_in[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input258_A wr_data[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1523__B1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input21_A core0_data_print[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1811__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0935__B _0951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output477_A _2145_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput407 _1731_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[31] sky130_fd_sc_hd__buf_2
Xoutput429 _1979_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[22] sky130_fd_sc_hd__buf_2
XANTENNA_output644_A _1090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1531_ _2097_/Q _1526_/X input55/X _1527_/X vssd1 vssd1 vccd1 vccd1 _2097_/D sky130_fd_sc_hd__a22o_1
Xoutput418 _1939_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[12] sky130_fd_sc_hd__buf_2
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1462_ input71/X _1459_/X _2048_/Q _1460_/X vssd1 vssd1 vccd1 vccd1 _2048_/D sky130_fd_sc_hd__o22a_1
XFILLER_4_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1393_ _2130_/Q _1389_/X input56/X _1390_/X vssd1 vssd1 vccd1 vccd1 _2130_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1514__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2014_ _2013_/X _2014_/A1 _2014_/S vssd1 vssd1 vccd1 vccd1 _2014_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1729_ _1729_/A vssd1 vssd1 vccd1 vccd1 _1729_/X sky130_fd_sc_hd__buf_2
XANTENNA__1692__A _1692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1505__B1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1808__A1 _1686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2091__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_135_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input69_A dout0_to_sram[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1806__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_110_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1107__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output594_A _1756_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0962_ _1732_/A _1720_/A vssd1 vssd1 vccd1 vccd1 _0963_/A sky130_fd_sc_hd__and2_1
XFILLER_32_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0893_ _0893_/A _0909_/B vssd1 vssd1 vccd1 vccd1 _0894_/A sky130_fd_sc_hd__and2_1
XFILLER_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1514_ _2084_/Q _1486_/A input76/X _1487_/A vssd1 vssd1 vccd1 vccd1 _2084_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1445_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1445_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1017__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1376_ _1390_/A vssd1 vssd1 vccd1 vccd1 _1376_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1687__A _1687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1577__684 vssd1 vssd1 vccd1 vccd1 _1577__684/HI la_data_out[25] sky130_fd_sc_hd__conb_1
XFILLER_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input123_A la_data_in[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output342_A _1682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1230_ _1232_/A _1230_/B vssd1 vssd1 vccd1 vccd1 _1242_/B sky130_fd_sc_hd__or2_1
XFILLER_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1161_ _1150_/A _1168_/A _1170_/B vssd1 vssd1 vccd1 vccd1 _1161_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1092_ _1092_/A vssd1 vssd1 vccd1 vccd1 _1092_/X sky130_fd_sc_hd__buf_2
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1994_ _1993_/X _1994_/A1 _2010_/S vssd1 vssd1 vccd1 vccd1 _1994_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0945_ _1732_/A _1716_/A vssd1 vssd1 vccd1 vccd1 _0946_/A sky130_fd_sc_hd__and2_1
XFILLER_119_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0876_ _0876_/A vssd1 vssd1 vccd1 vccd1 _0891_/A sky130_fd_sc_hd__inv_4
XFILLER_134_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1611__718 vssd1 vssd1 vccd1 vccd1 _1611__718/HI la_data_out[59] sky130_fd_sc_hd__conb_1
XFILLER_114_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1428_ input75/X _1422_/X _2024_/Q _1425_/X vssd1 vssd1 vccd1 vccd1 _2024_/D sky130_fd_sc_hd__o22a_1
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1359_ _1541_/A vssd1 vssd1 vccd1 vccd1 _1520_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1210__A _1210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput590 _1753_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[19] sky130_fd_sc_hd__buf_2
XANTENNA_input240_A wr_data[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1478__A2 _1470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0943__B _0951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1938__A0 _1937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1402__A2 _1396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output557_A _2102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1213_ _1221_/A _1218_/A _1213_/C _1213_/D vssd1 vssd1 vccd1 vccd1 _1225_/B sky130_fd_sc_hd__or4_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1144_ _1152_/A vssd1 vssd1 vccd1 vccd1 _1144_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1075_ _2019_/Q _1075_/B vssd1 vssd1 vccd1 vccd1 _1076_/A sky130_fd_sc_hd__and2_1
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1929__A0 _1928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2152__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1977_ _1976_/X _1977_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__mux2_1
X_0928_ _1732_/A _1712_/A vssd1 vssd1 vccd1 vccd1 _0929_/A sky130_fd_sc_hd__and2_1
XFILLER_134_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0859_ _0859_/A vssd1 vssd1 vccd1 vccd1 _0859_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1904__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput307 wr_data[98] vssd1 vssd1 vccd1 vccd1 _0887_/A sky130_fd_sc_hd__buf_4
XFILLER_130_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input190_A wr_data[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input288_A wr_data[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1633__740 vssd1 vssd1 vccd1 vccd1 _1633__740/HI la_data_out[81] sky130_fd_sc_hd__conb_1
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input51_A core0_data_print[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1814__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1115__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2025__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1900_ _0894_/X _1900_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1900_/X sky130_fd_sc_hd__mux2_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ _1830_/X input2/X _1938_/S vssd1 vssd1 vccd1 vccd1 _1831_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1387__A1 _2126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1762_ _1762_/A vssd1 vssd1 vccd1 vccd1 _1762_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1693_ _1693_/A vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1009__B _1009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1025__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0864__A _1700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1127_ _2019_/Q _1127_/B vssd1 vssd1 vccd1 vccd1 _1128_/A sky130_fd_sc_hd__and2_1
XANTENNA__1311__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1058_ _1058_/A vssd1 vssd1 vccd1 vccd1 _1058_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1695__A _1695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1378__A1 _2119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1617__724 vssd1 vssd1 vccd1 vccd1 _1617__724/HI la_data_out[65] sky130_fd_sc_hd__conb_1
XFILLER_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2048__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput115 la_data_in[48] vssd1 vssd1 vccd1 vccd1 _1716_/A sky130_fd_sc_hd__clkbuf_4
Xinput104 la_data_in[38] vssd1 vssd1 vccd1 vccd1 _1706_/A sky130_fd_sc_hd__buf_4
Xinput126 la_data_in[58] vssd1 vssd1 vccd1 vccd1 _1726_/A sky130_fd_sc_hd__clkbuf_4
Xinput148 la_data_in[78] vssd1 vssd1 vccd1 vccd1 _1748_/A sky130_fd_sc_hd__buf_4
Xinput137 la_data_in[68] vssd1 vssd1 vccd1 vccd1 _1738_/A sky130_fd_sc_hd__buf_4
Xinput159 la_data_in[88] vssd1 vssd1 vccd1 vccd1 _1758_/A sky130_fd_sc_hd__buf_6
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input203_A wr_data[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input99_A la_data_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1809__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1369__A1 _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_125_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0949__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output422_A _1955_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2030_ _2155_/CLK _2030_/D vssd1 vssd1 vccd1 vccd1 _2030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1814_ _1813_/X _1687_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1814_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1745_ _1745_/A vssd1 vssd1 vccd1 vccd1 _1745_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1532__A1 _2098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input153_A la_data_in[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1523__A1 _2091_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input14_A addr_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0951__B _0951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput408 _1703_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[3] sky130_fd_sc_hd__buf_2
XFILLER_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1530_ _2096_/Q _1526_/X input54/X _1527_/X vssd1 vssd1 vccd1 vccd1 _2096_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput419 _1943_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[13] sky130_fd_sc_hd__buf_2
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1461_ input70/X _1459_/X _2047_/Q _1460_/X vssd1 vssd1 vccd1 vccd1 _2047_/D sky130_fd_sc_hd__o22a_1
X_1392_ _2129_/Q _1389_/X input55/X _1390_/X vssd1 vssd1 vccd1 vccd1 _2129_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1514__A1 _2084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1514__B2 _1487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2013_ _2012_/X _2013_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _2013_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1450__B1 _2040_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1728_ _1728_/A vssd1 vssd1 vccd1 vccd1 _1728_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1505__A1 _2077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A addr_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1912__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1441__B1 _2033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input270_A wr_data[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1107__B _1107_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1822__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1123__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0962__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0961_ _0961_/A vssd1 vssd1 vccd1 vccd1 _0961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0892_ _1009_/B vssd1 vssd1 vccd1 vccd1 _0909_/B sky130_fd_sc_hd__buf_2
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1513_ _2083_/Q _1507_/X input74/X _1508_/X vssd1 vssd1 vccd1 vccd1 _2083_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2109__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1444_ input58/X _1438_/X _2036_/Q _1439_/X vssd1 vssd1 vccd1 vccd1 _2036_/D sky130_fd_sc_hd__o22a_1
XFILLER_68_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1017__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1375_ _1411_/A vssd1 vssd1 vccd1 vccd1 _1390_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1499__B1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1033__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1907__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A la_data_in[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1414__B1 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1965__A1 _1965_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input81_A dout0_to_sram[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1817__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1160_ _1160_/A _1175_/A vssd1 vssd1 vccd1 vccd1 _1170_/B sky130_fd_sc_hd__or2_1
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1091_ _2019_/Q _1091_/B vssd1 vssd1 vccd1 vccd1 _1092_/A sky130_fd_sc_hd__and2_1
XFILLER_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater652_A _1942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1993_ _1992_/X _1993_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1993_/X sky130_fd_sc_hd__mux2_1
X_0944_ _0944_/A vssd1 vssd1 vccd1 vccd1 _0944_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1405__B1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0875_ _0875_/A _2152_/Q _0875_/C vssd1 vssd1 vccd1 vccd1 _0876_/A sky130_fd_sc_hd__or3_4
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1650__757 vssd1 vssd1 vccd1 vccd1 _1650__757/HI la_data_out[98] sky130_fd_sc_hd__conb_1
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1427_ input64/X _1422_/X _2023_/Q _1425_/X vssd1 vssd1 vccd1 vccd1 _2023_/D sky130_fd_sc_hd__o22a_1
XANTENNA__2081__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1358_ _1540_/A vssd1 vssd1 vccd1 vccd1 _1541_/A sky130_fd_sc_hd__inv_2
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1289_ _1319_/A _1289_/B vssd1 vssd1 vccd1 vccd1 _1310_/A sky130_fd_sc_hd__or2_1
XANTENNA__1698__A _1698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput580 _1734_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[0] sky130_fd_sc_hd__buf_2
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput591 _1735_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[1] sky130_fd_sc_hd__buf_2
XFILLER_87_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input233_A wr_data[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1938__A1 _1938_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output452_A _2122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1212_ _1212_/A _1212_/B vssd1 vssd1 vccd1 vccd1 _1213_/C sky130_fd_sc_hd__or2_1
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1143_ input1/X vssd1 vssd1 vccd1 vccd1 _1152_/A sky130_fd_sc_hd__inv_2
XFILLER_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1074_ _1074_/A vssd1 vssd1 vccd1 vccd1 _1074_/X sky130_fd_sc_hd__buf_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1976_ _0973_/X _1976_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1976_/X sky130_fd_sc_hd__mux2_4
X_0927_ _0927_/A vssd1 vssd1 vccd1 vccd1 _0927_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0858_ _1733_/A _2151_/Q vssd1 vssd1 vccd1 vccd1 _0859_/A sky130_fd_sc_hd__and2_1
XFILLER_20_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput308 wr_data[99] vssd1 vssd1 vccd1 vccd1 _0893_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_130_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1920__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input183_A wr_data[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input44_A core0_data_print[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1115__B _1115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1830__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1131__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0970__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1830_ _1829_/X _1249_/Y _2013_/S vssd1 vssd1 vccd1 vccd1 _1830_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1761_ _1761_/A vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1692_ _1692_/A vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_98_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1025__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1126_ _1126_/A vssd1 vssd1 vccd1 vccd1 _1126_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0864__B _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1057_ _1733_/A _2151_/Q _1757_/A vssd1 vssd1 vccd1 vccd1 _1058_/A sky130_fd_sc_hd__and3_1
XFILLER_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1041__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1959_ _1958_/X _0950_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1959_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1656__763 vssd1 vssd1 vccd1 vccd1 _1656__763/HI la_data_out[105] sky130_fd_sc_hd__conb_1
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1915__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput127 la_data_in[59] vssd1 vssd1 vccd1 vccd1 _1727_/A sky130_fd_sc_hd__buf_2
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput116 la_data_in[49] vssd1 vssd1 vccd1 vccd1 _1717_/A sky130_fd_sc_hd__clkbuf_4
Xinput105 la_data_in[39] vssd1 vssd1 vccd1 vccd1 _1707_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput138 la_data_in[69] vssd1 vssd1 vccd1 vccd1 _1739_/A sky130_fd_sc_hd__buf_6
Xinput149 la_data_in[79] vssd1 vssd1 vccd1 vccd1 _1749_/A sky130_fd_sc_hd__buf_6
XFILLER_76_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_125_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1825__S _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0949__B _1717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2142__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output415_A _1891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1599__706 vssd1 vssd1 vccd1 vccd1 _1599__706/HI la_data_out[47] sky130_fd_sc_hd__conb_1
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1813_ _1812_/X _1210_/A _1938_/S vssd1 vssd1 vccd1 vccd1 _1813_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1744_ _1744_/A vssd1 vssd1 vccd1 vccd1 _1744_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1296__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2089_ _2149_/CLK _2089_/D vssd1 vssd1 vccd1 vccd1 _2089_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1109_ _2019_/Q _1109_/B vssd1 vssd1 vccd1 vccd1 _1110_/A sky130_fd_sc_hd__and2_1
XFILLER_54_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_135_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input146_A la_data_in[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output365_A _1056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput409 _1704_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[4] sky130_fd_sc_hd__buf_2
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1460_ _1460_/A vssd1 vssd1 vccd1 vccd1 _1460_/X sky130_fd_sc_hd__clkbuf_2
X_1391_ _2128_/Q _1389_/X input54/X _1390_/X vssd1 vssd1 vccd1 vccd1 _2128_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output532_A _2080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2012_ _1010_/X _2012_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__mux2_2
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2038__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1450__A1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1727_ _1727_/A vssd1 vssd1 vccd1 vccd1 _1727_/X sky130_fd_sc_hd__buf_2
XFILLER_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1441__A1 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input263_A wr_data[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1123__B _1123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1561__668 vssd1 vssd1 vccd1 vccd1 _1561__668/HI la_data_out[9] sky130_fd_sc_hd__conb_1
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0960_ _0960_/A _0972_/B vssd1 vssd1 vccd1 vccd1 _0961_/A sky130_fd_sc_hd__and2_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output482_A _2034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0891_ _0891_/A vssd1 vssd1 vccd1 vccd1 _1009_/B sky130_fd_sc_hd__buf_2
XFILLER_126_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1512_ _2082_/Q _1507_/X input73/X _1508_/X vssd1 vssd1 vccd1 vccd1 _2082_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1443_ input57/X _1438_/X _2035_/Q _1439_/X vssd1 vssd1 vccd1 vccd1 _2035_/D sky130_fd_sc_hd__o22a_1
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1374_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1411_/A sky130_fd_sc_hd__inv_2
XANTENNA__1499__A1 _2073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1017__C _1737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_56_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1033__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1923__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input109_A la_data_in[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1414__A1 _2145_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input74_A dout0_to_sram[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1833__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1090_ _1090_/A vssd1 vssd1 vccd1 vccd1 _1090_/X sky130_fd_sc_hd__buf_2
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1992_ _0990_/X _1992_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1992_/X sky130_fd_sc_hd__mux2_4
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1405__A1 _2138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0943_ _0943_/A _0951_/B vssd1 vssd1 vccd1 vccd1 _0944_/A sky130_fd_sc_hd__and2_1
XFILLER_118_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0874_ _0874_/A vssd1 vssd1 vccd1 vccd1 _2012_/S sky130_fd_sc_hd__buf_12
XFILLER_115_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0867__B _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1426_ input53/X _1422_/X _2022_/Q _1425_/X vssd1 vssd1 vccd1 vccd1 _2022_/D sky130_fd_sc_hd__o22a_1
X_1357_ _1519_/A vssd1 vssd1 vccd1 vccd1 _1357_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1892__A1 _1892_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1288_ input5/X _1275_/Y _1308_/A vssd1 vssd1 vccd1 vccd1 _1288_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0883__A _0883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1583__690 vssd1 vssd1 vccd1 vccd1 _1583__690/HI la_data_out[31] sky130_fd_sc_hd__conb_1
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1918__S _1934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput570 _2114_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[92] sky130_fd_sc_hd__buf_2
Xoutput581 _1744_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[10] sky130_fd_sc_hd__buf_2
Xoutput592 _1754_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[20] sky130_fd_sc_hd__buf_2
XFILLER_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input226_A wr_data[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1399__B1 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1828__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1129__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0968__A _0968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1211_ _1221_/B vssd1 vssd1 vccd1 vccd1 _1218_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1874__A1 _1697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1567__674 vssd1 vssd1 vccd1 vccd1 _1567__674/HI la_data_out[15] sky130_fd_sc_hd__conb_1
X_1142_ _0841_/X _0873_/C _1958_/S vssd1 vssd1 vccd1 vccd1 _1142_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1073_ _1733_/A _2151_/Q _1765_/A vssd1 vssd1 vccd1 vccd1 _1074_/A sky130_fd_sc_hd__and3_1
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1975_ _1974_/X _0967_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1975_/X sky130_fd_sc_hd__mux2_4
XFILLER_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0926_ _0926_/A _0930_/B vssd1 vssd1 vccd1 vccd1 _0927_/A sky130_fd_sc_hd__and2_1
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0857_ _0857_/A vssd1 vssd1 vccd1 vccd1 _0857_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1039__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput309 wr_data[9] vssd1 vssd1 vccd1 vccd1 _1926_/A1 sky130_fd_sc_hd__buf_2
X_1409_ _2142_/Q _1403_/X input69/X _1404_/X vssd1 vssd1 vccd1 vccd1 _2142_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input176_A req_out_core0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input37_A core0_data_print[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1856__A1 _1694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1131__B _1131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1601__708 vssd1 vssd1 vccd1 vccd1 _1601__708/HI la_data_out[49] sky130_fd_sc_hd__conb_1
XANTENNA__0970__B _1722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output395_A _1720_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1760_ _1760_/A vssd1 vssd1 vccd1 vccd1 _1760_/X sky130_fd_sc_hd__buf_4
XANTENNA__2071__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output562_A _2107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1792__A0 _1177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1691_ _1691_/A vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__buf_4
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1544__B1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1025__C _1741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1125_ _2019_/Q _1125_/B vssd1 vssd1 vccd1 vccd1 _1126_/A sky130_fd_sc_hd__and2_1
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1056_ _1056_/A vssd1 vssd1 vccd1 vccd1 _1056_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1041__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1958_ _1957_/X _1958_/A1 _1958_/S vssd1 vssd1 vccd1 vccd1 _1958_/X sky130_fd_sc_hd__mux2_2
XFILLER_31_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0909_ _0909_/A _0909_/B vssd1 vssd1 vccd1 vccd1 _0910_/A sky130_fd_sc_hd__and2_1
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1889_ _1888_/X _1889_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__mux2_2
XFILLER_134_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1535__B1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput117 la_data_in[4] vssd1 vssd1 vccd1 vccd1 _1684_/A sky130_fd_sc_hd__buf_4
XFILLER_130_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput106 la_data_in[3] vssd1 vssd1 vccd1 vccd1 _1683_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput128 la_data_in[5] vssd1 vssd1 vccd1 vccd1 _1685_/A sky130_fd_sc_hd__buf_6
Xinput139 la_data_in[6] vssd1 vssd1 vccd1 vccd1 _1686_/A sky130_fd_sc_hd__buf_2
XANTENNA__1931__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1838__A1 _1691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2094__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input293_A wr_data[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1774__A0 _1150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_137_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2002__S _2010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1841__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output310_A _1773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1679__786 vssd1 vssd1 vccd1 vccd1 _1679__786/HI spare_wen0_to_sram sky130_fd_sc_hd__conb_1
X_1812_ _1811_/X _1214_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1812_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1743_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1743_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1517__B1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0875__B _2152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2088_ _2149_/CLK _2088_/D vssd1 vssd1 vccd1 vccd1 _2088_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1108_ _1108_/A vssd1 vssd1 vccd1 vccd1 _1108_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1623__730 vssd1 vssd1 vccd1 vccd1 _1623__730/HI la_data_out[71] sky130_fd_sc_hd__conb_1
XANTENNA__0891__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1039_ _1733_/A _2151_/Q _1748_/A vssd1 vssd1 vccd1 vccd1 _1040_/A sky130_fd_sc_hd__and3_1
XFILLER_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1926__S _1958_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input139_A la_data_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input306_A wr_data[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1836__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1137__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output358_A _1044_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1390_ _1390_/A vssd1 vssd1 vccd1 vccd1 _1390_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output525_A _2073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2011_ _2010_/X _1004_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _2011_/X sky130_fd_sc_hd__mux2_4
X_1607__714 vssd1 vssd1 vccd1 vccd1 _1607__714/HI la_data_out[55] sky130_fd_sc_hd__conb_1
XFILLER_75_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1726_ _1726_/A vssd1 vssd1 vccd1 vccd1 _1726_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1047__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1910__A0 _1909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1977__A0 _1976_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2132__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input256_A wr_data[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1420__A _2021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0890_ _0890_/A vssd1 vssd1 vccd1 vccd1 _0890_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output475_A _2143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output642_A _1086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1511_ _2081_/Q _1507_/X input72/X _1508_/X vssd1 vssd1 vccd1 vccd1 _2081_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_126_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1442_ input56/X _1438_/X _2034_/Q _1439_/X vssd1 vssd1 vccd1 vccd1 _2034_/D sky130_fd_sc_hd__o22a_1
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1373_ _1389_/A vssd1 vssd1 vccd1 vccd1 _1373_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1033__C _1745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2155__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1959__A0 _1958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1709_ _1709_/A vssd1 vssd1 vccd1 vccd1 _1709_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_136_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input67_A dout0_to_sram[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2010__S _2010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2028__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1350__A1 _1349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1150__A _1150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output592_A _1754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1991_ _1990_/X _0984_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1991_/X sky130_fd_sc_hd__mux2_2
X_0942_ _0942_/A vssd1 vssd1 vccd1 vccd1 _0942_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0873_ _0875_/A _2152_/Q _0873_/C vssd1 vssd1 vccd1 vccd1 _0874_/A sky130_fd_sc_hd__and3_1
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1325__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1425_ _1439_/A vssd1 vssd1 vccd1 vccd1 _1425_/X sky130_fd_sc_hd__clkbuf_4
X_1356_ _1540_/A vssd1 vssd1 vccd1 vccd1 _1519_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1287_ _1319_/A _1319_/D vssd1 vssd1 vccd1 vccd1 _1308_/A sky130_fd_sc_hd__or2_1
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0883__B _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_133_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_105_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1934__S _1934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput560 _2105_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[83] sky130_fd_sc_hd__buf_2
Xoutput571 _2115_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[93] sky130_fd_sc_hd__buf_2
XFILLER_78_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput593 _1755_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[21] sky130_fd_sc_hd__buf_2
Xoutput582 _1745_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[11] sky130_fd_sc_hd__buf_2
XANTENNA__1235__A _1235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input121_A la_data_in[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input219_A wr_data[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1399__A1 _2134_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1399__B2 _1397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2005__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1844__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0968__B _0972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output340_A _1699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output438_A _2011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1210_ _1210_/A vssd1 vssd1 vccd1 vccd1 _1221_/B sky130_fd_sc_hd__inv_2
XFILLER_93_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1141_ _1732_/A vssd1 vssd1 vccd1 vccd1 _1141_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1072_ _1072_/A vssd1 vssd1 vccd1 vccd1 _1072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1974_ _1973_/X _1974_/A1 _1990_/S vssd1 vssd1 vccd1 vccd1 _1974_/X sky130_fd_sc_hd__mux2_2
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0925_ _0925_/A vssd1 vssd1 vccd1 vccd1 _0925_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0856_ _2016_/X _0856_/B vssd1 vssd1 vccd1 vccd1 _2151_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1039__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1408_ _2141_/Q _1403_/X input68/X _1404_/X vssd1 vssd1 vccd1 vccd1 _2141_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1055__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1339_ _1339_/A vssd1 vssd1 vccd1 vccd1 _1339_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1929__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_133_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input169_A la_data_in[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput390 _1716_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[16] sky130_fd_sc_hd__buf_2
XFILLER_75_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1640__747 vssd1 vssd1 vccd1 vccd1 _1640__747/HI la_data_out[88] sky130_fd_sc_hd__conb_1
XANTENNA__1839__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output388_A _1714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1690_ _1690_/A vssd1 vssd1 vccd1 vccd1 _1690_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output555_A _2101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0979__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1544__A1 _2106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1124_ _1124_/A vssd1 vssd1 vccd1 vccd1 _1124_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1055_ _1733_/A _2151_/Q _1756_/A vssd1 vssd1 vccd1 vccd1 _1056_/A sky130_fd_sc_hd__and3_1
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1041__C _1749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1957_ _1956_/X _1957_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1957_/X sky130_fd_sc_hd__mux2_2
XFILLER_135_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1888_ _0880_/X _1888_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1888_/X sky130_fd_sc_hd__mux2_2
X_0908_ _0908_/A vssd1 vssd1 vccd1 vccd1 _0908_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0889__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1535__B2 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput118 la_data_in[50] vssd1 vssd1 vccd1 vccd1 _1718_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput107 la_data_in[40] vssd1 vssd1 vccd1 vccd1 _1708_/A sky130_fd_sc_hd__buf_6
Xinput129 la_data_in[60] vssd1 vssd1 vccd1 vccd1 _1728_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_112_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input286_A wr_data[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0981__B _0993_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1462__B1 _2048_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1811_ _1810_/X _1217_/Y _2012_/S vssd1 vssd1 vccd1 vccd1 _1811_/X sky130_fd_sc_hd__mux2_1
X_1742_ _1742_/A vssd1 vssd1 vccd1 vccd1 _1742_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1517__A1 _2087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2087_ _1767_/X _2087_/D vssd1 vssd1 vccd1 vccd1 _2087_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1107_ _2019_/Q _1107_/B vssd1 vssd1 vccd1 vccd1 _1108_/A sky130_fd_sc_hd__and2_1
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1038_ _1038_/A vssd1 vssd1 vccd1 vccd1 _1038_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1942__S _1942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2061__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input201_A wr_data[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1444__B1 _2036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input97_A la_data_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2013__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1137__B _1137_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1852__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output420_A _1947_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2010_ _2009_/X _2010_/A1 _2010_/S vssd1 vssd1 vccd1 vccd1 _2010_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1646__753 vssd1 vssd1 vccd1 vccd1 _1646__753/HI la_data_out[94] sky130_fd_sc_hd__conb_1
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1435__B1 _2029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1725_ _1725_/A vssd1 vssd1 vccd1 vccd1 _1725_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1047__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2084__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1063__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ _2149_/CLK _2139_/D vssd1 vssd1 vccd1 vccd1 _2139_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1977__A1 _1977_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1937__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_135_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input151_A la_data_in[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input249_A wr_data[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input12_A addr_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1420__B _2020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1417__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2008__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1847__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output468_A _2137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1510_ _2080_/Q _1507_/X input71/X _1508_/X vssd1 vssd1 vccd1 vccd1 _2080_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1441_ input55/X _1438_/X _2033_/Q _1439_/X vssd1 vssd1 vccd1 vccd1 _2033_/D sky130_fd_sc_hd__o22a_1
XANTENNA__0987__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output635_A _1132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1372_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1389_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput290 wr_data[82] vssd1 vssd1 vccd1 vccd1 _1960_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1408__B1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1959__A1 _0950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_133_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1708_ _1708_/A vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0897__A _0897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input4_A addr_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1895__A0 _1894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input199_A wr_data[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1431__A _1438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1990_ _1989_/X _1990_/A1 _1990_/S vssd1 vssd1 vccd1 vccd1 _1990_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ _1732_/A _1715_/A vssd1 vssd1 vccd1 vccd1 _0942_/A sky130_fd_sc_hd__and2_1
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1810__A0 _1210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0872_ _0872_/A vssd1 vssd1 vccd1 vccd1 _2013_/S sky130_fd_sc_hd__buf_12
XFILLER_115_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1424_ _1460_/A vssd1 vssd1 vccd1 vccd1 _1439_/A sky130_fd_sc_hd__buf_4
XFILLER_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1355_ _1371_/A _2020_/Q vssd1 vssd1 vccd1 vccd1 _1540_/A sky130_fd_sc_hd__or2_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_110_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2122__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1286_ _1319_/A _1284_/B _1285_/Y vssd1 vssd1 vccd1 vccd1 _1286_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_105_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput572 _2116_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[94] sky130_fd_sc_hd__buf_2
Xoutput550 _2096_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[74] sky130_fd_sc_hd__buf_2
XFILLER_132_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput561 _2106_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[84] sky130_fd_sc_hd__buf_2
XFILLER_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput594 _1756_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[22] sky130_fd_sc_hd__buf_2
X_1551__658 vssd1 vssd1 vccd1 vccd1 _1551__658/HI csb0_to_sram sky130_fd_sc_hd__conb_1
Xoutput583 _1746_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[12] sky130_fd_sc_hd__buf_2
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1950__S _2010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input114_A la_data_in[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1399__A2 _1396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_136_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output333_A _1692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2145__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1140_ _1140_/A vssd1 vssd1 vccd1 vccd1 _1419_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1860__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1071_ _1733_/A _2151_/Q _1764_/A vssd1 vssd1 vccd1 vccd1 _1072_/A sky130_fd_sc_hd__and3_1
XANTENNA_output500_A _2051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater650_A _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1973_ _1972_/X _1973_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1973_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0924_ _1732_/A _1711_/A vssd1 vssd1 vccd1 vccd1 _0925_/A sky130_fd_sc_hd__and2_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0855_ _0854_/Y _2151_/Q _0857_/A _2150_/Q vssd1 vssd1 vccd1 vccd1 _0856_/B sky130_fd_sc_hd__a22oi_1
XFILLER_134_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1039__C _1748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1336__A _1336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1407_ _2140_/Q _1403_/X input67/X _1404_/X vssd1 vssd1 vccd1 vccd1 _2140_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1055__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1770__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1338_ _1341_/A _1338_/B vssd1 vssd1 vccd1 vccd1 _1339_/A sky130_fd_sc_hd__or2_1
XFILLER_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1071__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1269_ _1274_/A _1269_/B vssd1 vssd1 vccd1 vccd1 _1282_/B sky130_fd_sc_hd__or2_1
XFILLER_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__2018__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1945__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1246__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput380 _1026_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[7] sky130_fd_sc_hd__buf_2
Xoutput391 _1717_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[17] sky130_fd_sc_hd__buf_2
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input231_A wr_data[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2016__S _2016_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1855__S _1942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0979__B _1724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1573__680 vssd1 vssd1 vccd1 vccd1 _1573__680/HI la_data_out[21] sky130_fd_sc_hd__conb_1
XANTENNA_output450_A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output548_A _2094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0995__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1123_ _2019_/Q _1123_/B vssd1 vssd1 vccd1 vccd1 _1124_/A sky130_fd_sc_hd__and2_1
XFILLER_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1054_ _1054_/A vssd1 vssd1 vccd1 vccd1 _1054_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1956_ _0952_/X _1956_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1956_/X sky130_fd_sc_hd__mux2_8
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0907_ _1732_/A _1707_/A vssd1 vssd1 vccd1 vccd1 _0908_/A sky130_fd_sc_hd__and2_1
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1887_ _1353_/X _1886_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1887_/X sky130_fd_sc_hd__mux2_2
XANTENNA__0889__B _1703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1535__A2 _1533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput108 la_data_in[41] vssd1 vssd1 vccd1 vccd1 _1709_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput119 la_data_in[51] vssd1 vssd1 vccd1 vccd1 _1719_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1557__664 vssd1 vssd1 vccd1 vccd1 _1557__664/HI la_data_out[5] sky130_fd_sc_hd__conb_1
XANTENNA_input279_A wr_data[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input181_A we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_137_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input42_A core0_data_print[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1704__A _1704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1462__A1 input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output498_A _2049_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1810_ _1210_/A _1220_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1810_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1214__A1 _1210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1741_ _1741_/A vssd1 vssd1 vccd1 vccd1 _1741_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2155_/CLK _2155_/D vssd1 vssd1 vccd1 vccd1 _2155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1106_ _1106_/A vssd1 vssd1 vccd1 vccd1 _1106_/X sky130_fd_sc_hd__clkbuf_4
X_2086_ _2149_/CLK _2086_/D vssd1 vssd1 vccd1 vccd1 _2086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1037_ _1733_/A _2151_/Q _1747_/A vssd1 vssd1 vccd1 vccd1 _1038_/A sky130_fd_sc_hd__and3_1
XFILLER_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1939_ _1938_/X _0929_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1939_/X sky130_fd_sc_hd__mux2_1
Xinput90 la_data_in[14] vssd1 vssd1 vccd1 vccd1 _1694_/A sky130_fd_sc_hd__buf_4
XFILLER_135_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1444__A1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_122_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1380__B1 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1435__A1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1724_ _1724_/A vssd1 vssd1 vccd1 vccd1 _1724_/X sky130_fd_sc_hd__buf_4
XFILLER_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1047__C _1752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1063__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2138_ _1767_/X _2138_/D vssd1 vssd1 vccd1 vccd1 _2138_/Q sky130_fd_sc_hd__dfxtp_4
X_2069_ _2149_/CLK _2069_/D vssd1 vssd1 vccd1 vccd1 _2069_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1426__A1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1426__B2 _1425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1953__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input144_A la_data_in[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1362__B1 input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1669__776 vssd1 vssd1 vccd1 vccd1 _1669__776/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XFILLER_94_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1417__A1 _2148_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output363_A _1052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1863__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1613__720 vssd1 vssd1 vccd1 vccd1 _1613__720/HI la_data_out[61] sky130_fd_sc_hd__conb_1
X_1440_ input54/X _1438_/X _2032_/Q _1439_/X vssd1 vssd1 vccd1 vccd1 _2032_/D sky130_fd_sc_hd__o22a_1
XANTENNA__0987__B _1726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1371_ _1371_/A _1468_/B vssd1 vssd1 vccd1 vccd1 _1410_/A sky130_fd_sc_hd__or2_2
XANTENNA_output530_A _2078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output628_A _1118_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_110_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput280 wr_data[73] vssd1 vssd1 vccd1 vccd1 _1924_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput291 wr_data[83] vssd1 vssd1 vccd1 vccd1 _1964_/A1 sky130_fd_sc_hd__buf_2
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1408__A1 _2141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2051__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1707_ _1707_/A vssd1 vssd1 vccd1 vccd1 _1707_/X sky130_fd_sc_hd__buf_2
XANTENNA__1773__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0897__B _0909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1948__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_135_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input261_A wr_data[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1886__A1 _1699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1712__A _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1858__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ _0940_/A vssd1 vssd1 vccd1 vccd1 _0940_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2074__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output480_A _2148_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0871_ _2154_/Q _2152_/Q _0873_/C vssd1 vssd1 vccd1 vccd1 _0872_/A sky130_fd_sc_hd__and3_1
XFILLER_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1423_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1460_/A sky130_fd_sc_hd__inv_2
XFILLER_122_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1354_ _2021_/Q vssd1 vssd1 vccd1 vccd1 _1371_/A sky130_fd_sc_hd__inv_2
XFILLER_110_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1285_ _1295_/B vssd1 vssd1 vccd1 vccd1 _1285_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1768__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1069__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1801__A1 _1189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1590__697 vssd1 vssd1 vccd1 vccd1 _1590__697/HI la_data_out[38] sky130_fd_sc_hd__conb_1
Xoutput562 _2107_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[85] sky130_fd_sc_hd__buf_2
XFILLER_105_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput551 _2097_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[75] sky130_fd_sc_hd__buf_2
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput540 _2087_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[65] sky130_fd_sc_hd__buf_2
Xoutput595 _1757_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[23] sky130_fd_sc_hd__buf_2
Xoutput573 _2117_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[95] sky130_fd_sc_hd__buf_2
XFILLER_115_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput584 _1747_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[13] sky130_fd_sc_hd__buf_2
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1868__A1 _1696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2097__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input107_A la_data_in[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input72_A dout0_to_sram[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1070_ _1070_/A vssd1 vssd1 vccd1 vccd1 _1070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1972_ _0969_/X _1972_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1972_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0923_ _0923_/A vssd1 vssd1 vccd1 vccd1 _0923_/X sky130_fd_sc_hd__clkbuf_1
X_0854_ _1733_/A vssd1 vssd1 vccd1 vccd1 _0854_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1547__B1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1406_ _2139_/Q _1403_/X input66/X _1404_/X vssd1 vssd1 vccd1 vccd1 _2139_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1055__C _1756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1337_ _1346_/A vssd1 vssd1 vccd1 vccd1 _1341_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1071__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1268_ _1277_/A vssd1 vssd1 vccd1 vccd1 _1274_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1199_ _1189_/A _1187_/Y _1221_/C vssd1 vssd1 vccd1 vccd1 _1199_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1538__B1 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1961__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput370 _1066_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[27] sky130_fd_sc_hd__buf_2
Xoutput392 _1718_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[18] sky130_fd_sc_hd__buf_2
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput381 _1028_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[8] sky130_fd_sc_hd__buf_2
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input224_A wr_data[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1529__B1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2112__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output443_A _1915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1871__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0995__B _1728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1122_ _1122_/A vssd1 vssd1 vccd1 vccd1 _1122_/X sky130_fd_sc_hd__clkbuf_4
X_1053_ _1733_/A _2151_/Q _1755_/A vssd1 vssd1 vccd1 vccd1 _1054_/A sky130_fd_sc_hd__and3_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2009__A1 _2009_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1955_ _1954_/X _0946_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1955_/X sky130_fd_sc_hd__mux2_2
XFILLER_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0906_ _0906_/A vssd1 vssd1 vccd1 vccd1 _0906_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1886_ _1885_/X _1699_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1886_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1781__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput109 la_data_in[42] vssd1 vssd1 vccd1 vccd1 _1710_/A sky130_fd_sc_hd__buf_6
XFILLER_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1956__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2135__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1257__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input174_A la_oenb[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_134_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input35_A core0_data_print[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output393_A _1719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1866__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1740_ _1740_/A vssd1 vssd1 vccd1 vccd1 _1740_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output560_A _2105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1922__A0 _1921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2154_ _2155_/CLK _2154_/D vssd1 vssd1 vccd1 vccd1 _2154_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1105_ _2019_/Q _1105_/B vssd1 vssd1 vccd1 vccd1 _1106_/A sky130_fd_sc_hd__and2_1
X_2085_ _2149_/CLK _2085_/D vssd1 vssd1 vccd1 vccd1 _2085_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1036_ _1036_/A vssd1 vssd1 vccd1 vccd1 _1036_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1989__A0 _1988_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1776__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1938_ _1937_/X _1938_/A1 _1938_/S vssd1 vssd1 vccd1 vccd1 _1938_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1077__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1869_ _1324_/Y _1868_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1869_/X sky130_fd_sc_hd__mux2_2
Xinput91 la_data_in[15] vssd1 vssd1 vccd1 vccd1 _1695_/A sky130_fd_sc_hd__buf_4
Xinput80 dout0_to_sram[5] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__buf_12
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1630__737 vssd1 vssd1 vccd1 vccd1 _1630__737/HI la_data_out[78] sky130_fd_sc_hd__conb_1
XFILLER_89_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1913__A0 _1912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input291_A wr_data[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1715__A _1715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1380__A1 _2121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output406_A _1730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1199__A1 _1189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1723_ _1723_/A vssd1 vssd1 vccd1 vccd1 _1723_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1063__C _1760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2137_ _1767_/X _2137_/D vssd1 vssd1 vccd1 vccd1 _2137_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2068_ _1767_/X _2068_/D vssd1 vssd1 vccd1 vccd1 _2068_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1019_ _1733_/A _2151_/Q _1738_/A vssd1 vssd1 vccd1 vccd1 _1020_/A sky130_fd_sc_hd__and3_1
XANTENNA__1426__A2 _1422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1362__A1 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input137_A la_data_in[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input304_A wr_data[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1370_ _2020_/Q vssd1 vssd1 vccd1 vccd1 _1468_/B sky130_fd_sc_hd__inv_2
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1353__A1 _1349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output523_A _2026_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput281 wr_data[74] vssd1 vssd1 vccd1 vccd1 _1928_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput270 wr_data[64] vssd1 vssd1 vccd1 vccd1 _1888_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput292 wr_data[84] vssd1 vssd1 vccd1 vccd1 _1968_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1706_ _1706_/A vssd1 vssd1 vccd1 vccd1 _1706_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1499_ _2073_/Q _1493_/X input63/X _1494_/X vssd1 vssd1 vccd1 vccd1 _2073_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1595__702 vssd1 vssd1 vccd1 vccd1 _1595__702/HI la_data_out[43] sky130_fd_sc_hd__conb_1
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1964__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1636__743 vssd1 vssd1 vccd1 vccd1 _1636__743/HI la_data_out[84] sky130_fd_sc_hd__conb_1
XFILLER_136_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_124_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_135_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input254_A wr_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1335__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0870_ _0870_/A _0870_/B _2153_/Q vssd1 vssd1 vccd1 vccd1 _1958_/S sky130_fd_sc_hd__nor3_4
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output473_A _2033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1874__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output640_A _1082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1422_ _1438_/A vssd1 vssd1 vccd1 vccd1 _1422_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1353_ _1349_/A _1347_/Y _1349_/Y _1347_/A vssd1 vssd1 vccd1 vccd1 _1353_/X sky130_fd_sc_hd__o22a_1
XFILLER_110_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1284_ _1284_/A _1284_/B vssd1 vssd1 vccd1 vccd1 _1295_/B sky130_fd_sc_hd__or2_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1069__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0999_ _1732_/A _1729_/A vssd1 vssd1 vccd1 vccd1 _1000_/A sky130_fd_sc_hd__and2_1
XFILLER_118_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1784__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput552 _2098_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[76] sky130_fd_sc_hd__buf_2
XFILLER_133_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput563 _2108_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[86] sky130_fd_sc_hd__buf_2
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput541 _2088_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[66] sky130_fd_sc_hd__buf_2
XFILLER_59_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1085__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput530 _2078_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[56] sky130_fd_sc_hd__buf_2
Xoutput574 _2118_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[96] sky130_fd_sc_hd__buf_2
Xoutput596 _1758_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[24] sky130_fd_sc_hd__buf_2
Xoutput585 _1748_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[14] sky130_fd_sc_hd__buf_2
XFILLER_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_131_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1959__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_6_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_136_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input65_A dout0_to_sram[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1723__A _1723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2041__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output319_A _1881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1869__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1492__B1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output590_A _1753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1971_ _1970_/X _0963_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1971_/X sky130_fd_sc_hd__mux2_2
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0922_ _0922_/A _0930_/B vssd1 vssd1 vccd1 vccd1 _0923_/A sky130_fd_sc_hd__and2_1
XANTENNA__1795__A1 _1177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0853_ _0853_/A vssd1 vssd1 vccd1 vccd1 _2152_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1547__A1 _2109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1405_ _2138_/Q _1403_/X input65/X _1404_/X vssd1 vssd1 vccd1 vccd1 _2138_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1336_ _1336_/A vssd1 vssd1 vccd1 vccd1 _1346_/A sky130_fd_sc_hd__inv_2
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput1 addr_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_84_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1267_ input4/X vssd1 vssd1 vccd1 vccd1 _1277_/A sky130_fd_sc_hd__inv_2
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1071__C _1764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1779__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1198_ _1212_/B _1198_/B vssd1 vssd1 vccd1 vccd1 _1221_/C sky130_fd_sc_hd__or2_1
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1483__B1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1538__B2 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1538__A1 _2102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput371 _1068_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[28] sky130_fd_sc_hd__buf_2
Xoutput360 _1048_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[18] sky130_fd_sc_hd__buf_2
XFILLER_121_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput382 _1030_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[9] sky130_fd_sc_hd__buf_2
Xoutput393 _1719_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[19] sky130_fd_sc_hd__buf_2
XFILLER_87_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2064__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input217_A wr_data[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1474__B1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1777__A1 _1150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1529__A1 _2095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output603_A _1764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1121_ _2019_/Q _1121_/B vssd1 vssd1 vccd1 vccd1 _1122_/A sky130_fd_sc_hd__and2_1
XFILLER_81_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1052_ _1052_/A vssd1 vssd1 vccd1 vccd1 _1052_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1465__B1 _2051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1954_ _1953_/X _1954_/A1 _1954_/S vssd1 vssd1 vccd1 vccd1 _1954_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0905_ _0905_/A _0909_/B vssd1 vssd1 vccd1 vccd1 _0906_/A sky130_fd_sc_hd__and2_1
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_135_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1885_ _1884_/X _1349_/A _1954_/S vssd1 vssd1 vccd1 vccd1 _1885_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2087__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1940__A1 _1940_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1319_ _1319_/A _1319_/B _1319_/C _1319_/D vssd1 vssd1 vccd1 vccd1 _1343_/C sky130_fd_sc_hd__or4_2
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1456__B1 _2044_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1972__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_134_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input167_A la_data_in[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input28_A core0_data_print[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1447__B1 _2037_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1882__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1922__A1 _1922_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2153_ _2155_/CLK _2153_/D vssd1 vssd1 vccd1 vccd1 _2153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1104_ _1104_/A vssd1 vssd1 vccd1 vccd1 _1104_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2084_ _2149_/CLK _2084_/D vssd1 vssd1 vccd1 vccd1 _2084_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1035_ _1733_/A _2151_/Q _1746_/A vssd1 vssd1 vccd1 vccd1 _1036_/A sky130_fd_sc_hd__and3_1
XANTENNA__1989__A1 _1989_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1937_ _1936_/X _1937_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1937_/X sky130_fd_sc_hd__mux2_2
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1868_ _1867_/X _1696_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1868_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1077__B _1077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput70 dout0_to_sram[25] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_6
Xinput81 dout0_to_sram[6] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_6
XANTENNA__1792__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput92 la_data_in[16] vssd1 vssd1 vccd1 vccd1 _1696_/A sky130_fd_sc_hd__buf_4
X_1799_ _1798_/X _1194_/Y _2012_/S vssd1 vssd1 vccd1 vccd1 _1799_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1093__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2102__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1563__670 vssd1 vssd1 vccd1 vccd1 _1563__670/HI la_data_out[11] sky130_fd_sc_hd__conb_1
XFILLER_12_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1967__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_138_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input284_A wr_data[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1904__A1 _1904_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1731__A _1731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1840__A0 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1877__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1722_ _1722_/A vssd1 vssd1 vccd1 vccd1 _1722_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2125__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2136_ _1767_/X _2136_/D vssd1 vssd1 vccd1 vccd1 _2136_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2067_ _1767_/X _2067_/D vssd1 vssd1 vccd1 vccd1 _2067_/Q sky130_fd_sc_hd__dfxtp_1
X_1018_ _1018_/A vssd1 vssd1 vccd1 vccd1 _1018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1787__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1898__A0 _1897_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1822__A0 _1235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input95_A la_data_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1726__A _1726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1889__A0 _1888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2148__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output349_A _1689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput271 wr_data[65] vssd1 vssd1 vccd1 vccd1 _1892_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput260 wr_data[55] vssd1 vssd1 vccd1 vccd1 _1981_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput293 wr_data[85] vssd1 vssd1 vccd1 vccd1 _1972_/A1 sky130_fd_sc_hd__buf_6
Xinput282 wr_data[75] vssd1 vssd1 vccd1 vccd1 _1932_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1705_ _1705_/A vssd1 vssd1 vccd1 vccd1 _1705_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1355__B _2020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1498_ _2072_/Q _1493_/X input62/X _1494_/X vssd1 vssd1 vccd1 vccd1 _2072_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ _2149_/CLK _2119_/D vssd1 vssd1 vccd1 vccd1 _2119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1675__782 vssd1 vssd1 vccd1 vccd1 _1675__782/HI la_data_out[124] sky130_fd_sc_hd__conb_1
XFILLER_129_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1980__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input247_A wr_data[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input10_A addr_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output466_A _2135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1421_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1438_/A sky130_fd_sc_hd__buf_4
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1890__S _1934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1352_ _1349_/A _1344_/Y _1349_/Y _1344_/A vssd1 vssd1 vccd1 vccd1 _1352_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1283_ input5/X _1270_/Y _1303_/A vssd1 vssd1 vccd1 vccd1 _1283_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1069__C _1763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1659__766 vssd1 vssd1 vccd1 vccd1 _1659__766/HI la_data_out[108] sky130_fd_sc_hd__conb_1
XFILLER_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0998_ _0998_/A vssd1 vssd1 vccd1 vccd1 _0998_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput520 _2069_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[47] sky130_fd_sc_hd__buf_2
XFILLER_133_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_117_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput553 _2099_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[77] sky130_fd_sc_hd__buf_2
Xoutput542 _2089_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[67] sky130_fd_sc_hd__buf_2
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1085__B _1085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput531 _2079_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[57] sky130_fd_sc_hd__buf_2
Xoutput575 _2119_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[97] sky130_fd_sc_hd__buf_2
Xoutput564 _2109_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[87] sky130_fd_sc_hd__buf_2
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput586 _1749_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[15] sky130_fd_sc_hd__buf_2
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput597 _1759_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[25] sky130_fd_sc_hd__buf_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input2_A addr_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1603__710 vssd1 vssd1 vccd1 vccd1 _1603__710/HI la_data_out[51] sky130_fd_sc_hd__conb_1
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1975__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input197_A wr_data[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input58_A dout0_to_sram[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_112_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1492__A1 _2068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1970_ _1969_/X _1970_/A1 _2014_/S vssd1 vssd1 vccd1 vccd1 _1970_/X sky130_fd_sc_hd__mux2_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0921_ _0921_/A vssd1 vssd1 vccd1 vccd1 _0921_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1885__S _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output583_A _1746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0852_ _0851_/X _0852_/B vssd1 vssd1 vccd1 vccd1 _0853_/A sky130_fd_sc_hd__and2b_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1404_ _1411_/A vssd1 vssd1 vccd1 vccd1 _1404_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1335_ input9/X _1323_/Y _1346_/B vssd1 vssd1 vccd1 vccd1 _1335_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 addr_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1266_ input3/X _1255_/Y _1277_/B vssd1 vssd1 vccd1 vccd1 _1266_/X sky130_fd_sc_hd__o21a_1
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1197_ _1195_/A _1195_/B _1196_/Y vssd1 vssd1 vccd1 vccd1 _1197_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1483__A1 _2061_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1795__S _1922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1538__A2 _1533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput361 _1050_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[19] sky130_fd_sc_hd__buf_2
Xoutput350 _2155_/CLK vssd1 vssd1 vccd1 vccd1 clk sky130_fd_sc_hd__buf_2
Xoutput372 _1070_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[29] sky130_fd_sc_hd__buf_2
XFILLER_114_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput394 _1701_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[1] sky130_fd_sc_hd__buf_2
Xoutput383 _1700_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[0] sky130_fd_sc_hd__buf_2
XFILLER_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input112_A la_data_in[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1474__B2 _1473_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0903__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output429_A _1979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1120_ _1120_/A vssd1 vssd1 vccd1 vccd1 _1120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1051_ _1733_/A _2151_/Q _1754_/A vssd1 vssd1 vccd1 vccd1 _1052_/A sky130_fd_sc_hd__and3_1
XFILLER_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1465__A1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580__687 vssd1 vssd1 vccd1 vccd1 _1580__687/HI la_data_out[28] sky130_fd_sc_hd__conb_1
XFILLER_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1953_ _1952_/X _1953_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1953_/X sky130_fd_sc_hd__mux2_2
X_0904_ _0904_/A vssd1 vssd1 vccd1 vccd1 _0904_/X sky130_fd_sc_hd__clkbuf_1
X_1884_ _1883_/X _1350_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1884_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_110_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1318_ input8/X _1306_/Y _1329_/B vssd1 vssd1 vccd1 vccd1 _1318_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1249_ _1252_/A _1258_/C _1248_/Y vssd1 vssd1 vccd1 vccd1 _1249_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1456__A1 input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1456__B2 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_119_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2031__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1392__B1 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1447__A1 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1729__A _1729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output379_A _1024_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output546_A _2092_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2152_ _2155_/CLK _2152_/D vssd1 vssd1 vccd1 vccd1 _2152_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2083_ _2149_/CLK _2083_/D vssd1 vssd1 vccd1 vccd1 _2083_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1103_ _2019_/Q _1103_/B vssd1 vssd1 vccd1 vccd1 _1104_/A sky130_fd_sc_hd__and2_1
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1034_ _1034_/A vssd1 vssd1 vccd1 vccd1 _1034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1936_ _0931_/X _1936_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1936_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2054__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1867_ _1866_/X input8/X _1954_/S vssd1 vssd1 vccd1 vccd1 _1867_/X sky130_fd_sc_hd__mux2_1
Xinput60 dout0_to_sram[16] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_6
Xinput71 dout0_to_sram[26] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_6
Xinput82 dout0_to_sram[7] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__buf_6
X_1798_ _1189_/A _1197_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1798_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput93 la_data_in[17] vssd1 vssd1 vccd1 vccd1 _1697_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1093__B _1093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xrepeater650 _1954_/S vssd1 vssd1 vccd1 vccd1 _1990_/S sky130_fd_sc_hd__buf_4
XFILLER_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1429__A1 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1429__B2 _1425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1983__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input277_A wr_data[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_106_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1365__B1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input40_A core0_data_print[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2077__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output496_A _2047_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1721_ _1721_/A vssd1 vssd1 vccd1 vccd1 _1721_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1893__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2135_ _1767_/X _2135_/D vssd1 vssd1 vccd1 vccd1 _2135_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1586__693 vssd1 vssd1 vccd1 vccd1 _1586__693/HI la_data_out[34] sky130_fd_sc_hd__conb_1
XFILLER_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2066_ _1767_/X _2066_/D vssd1 vssd1 vccd1 vccd1 _2066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1017_ _1733_/A _2151_/Q _1737_/A vssd1 vssd1 vccd1 vccd1 _1018_/A sky130_fd_sc_hd__and3_1
XFILLER_35_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1831__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1919_ _1918_/X _0908_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1919_/X sky130_fd_sc_hd__mux2_4
XFILLER_135_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1898__A1 _1898_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1978__S _2014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input88_A la_data_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0911__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1889__A1 _1889_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1742__A _1742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput272 wr_data[66] vssd1 vssd1 vccd1 vccd1 _1896_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput261 wr_data[56] vssd1 vssd1 vccd1 vccd1 _1985_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput250 wr_data[46] vssd1 vssd1 vccd1 vccd1 _1945_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput294 wr_data[86] vssd1 vssd1 vccd1 vccd1 _1976_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput283 wr_data[76] vssd1 vssd1 vccd1 vccd1 _1936_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__1510__B1 input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output509_A _2059_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1888__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1620__727 vssd1 vssd1 vccd1 vccd1 _1620__727/HI la_data_out[68] sky130_fd_sc_hd__conb_1
XANTENNA__1189__A _1189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1813__A1 _1210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1704_ _1704_/A vssd1 vssd1 vccd1 vccd1 _1704_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1497_ _2071_/Q _1493_/X input61/X _1494_/X vssd1 vssd1 vccd1 vccd1 _2071_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2118_ _2149_/CLK _2118_/D vssd1 vssd1 vccd1 vccd1 _2118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0855__A2 _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2049_ _2155_/CLK _2049_/D vssd1 vssd1 vccd1 vccd1 _2049_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1798__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1099__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_136_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input142_A la_data_in[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2115__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1737__A _1737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output361_A _1050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1420_ _2021_/Q _2020_/Q vssd1 vssd1 vccd1 vccd1 _1459_/A sky130_fd_sc_hd__or2_2
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1351_ _1336_/A _1330_/Y _1349_/Y _1349_/A _1341_/X vssd1 vssd1 vccd1 vccd1 _1351_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output626_A _1078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1282_ _1319_/A _1282_/B vssd1 vssd1 vccd1 vccd1 _1303_/A sky130_fd_sc_hd__or2_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1798__A0 _1189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0997_ _0997_/A _1009_/B vssd1 vssd1 vccd1 vccd1 _0998_/A sky130_fd_sc_hd__and2_1
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput510 _2060_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[38] sky130_fd_sc_hd__buf_2
Xoutput554 _2100_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[78] sky130_fd_sc_hd__buf_2
XFILLER_133_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1970__A0 _1969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput543 _2090_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[68] sky130_fd_sc_hd__buf_2
Xoutput521 _2070_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[48] sky130_fd_sc_hd__buf_2
Xoutput532 _2080_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[58] sky130_fd_sc_hd__buf_2
Xoutput587 _1750_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[16] sky130_fd_sc_hd__buf_2
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput565 _2110_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[88] sky130_fd_sc_hd__buf_2
Xoutput576 _2120_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[98] sky130_fd_sc_hd__buf_2
XFILLER_101_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput598 _1760_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[26] sky130_fd_sc_hd__buf_2
X_1549_ _0867_/A _2017_/S _0841_/X vssd1 vssd1 vccd1 vccd1 _1549_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2138__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1991__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ _1732_/A _1710_/A vssd1 vssd1 vccd1 vccd1 _0921_/A sky130_fd_sc_hd__and2_1
X_0851_ _0875_/A _0849_/Y _0870_/B _0873_/C vssd1 vssd1 vccd1 vccd1 _0851_/X sky130_fd_sc_hd__o22a_1
XANTENNA_output576_A _2120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1403_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1403_/X sky130_fd_sc_hd__clkbuf_2
X_1334_ _1334_/A _1334_/B vssd1 vssd1 vccd1 vccd1 _1346_/B sky130_fd_sc_hd__or2_1
XFILLER_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1265_ _1265_/A _1265_/B vssd1 vssd1 vccd1 vccd1 _1277_/B sky130_fd_sc_hd__or2_1
XFILLER_110_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput3 addr_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_4
X_1626__733 vssd1 vssd1 vccd1 vccd1 _1626__733/HI la_data_out[74] sky130_fd_sc_hd__conb_1
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1196_ _1206_/B vssd1 vssd1 vccd1 vccd1 _1196_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput340 _1699_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[19] sky130_fd_sc_hd__buf_2
Xoutput362 _1014_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[1] sky130_fd_sc_hd__buf_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput351 _1012_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[0] sky130_fd_sc_hd__buf_2
XFILLER_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput395 _1720_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[20] sky130_fd_sc_hd__buf_2
Xoutput373 _1016_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[2] sky130_fd_sc_hd__buf_2
Xoutput384 _1710_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[10] sky130_fd_sc_hd__buf_2
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1474__A2 _1470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input105_A la_data_in[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1986__S _1990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0903__B _1706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input70_A dout0_to_sram[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1934__A0 _1933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_112_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1750__A _1750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output324_A _1797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1050_ _1050_/A vssd1 vssd1 vccd1 vccd1 _1050_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1896__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ _0948_/X _1952_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1952_/X sky130_fd_sc_hd__mux2_4
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0903_ _1732_/A _1706_/A vssd1 vssd1 vccd1 vccd1 _0904_/A sky130_fd_sc_hd__and2_1
X_1883_ _1882_/X _1351_/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1883_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1317_ _1319_/C _1317_/B vssd1 vssd1 vccd1 vccd1 _1329_/B sky130_fd_sc_hd__or2_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1248_ _1252_/A _1258_/C vssd1 vssd1 vccd1 vccd1 _1248_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1456__A2 _1452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1179_ _1179_/A vssd1 vssd1 vccd1 vccd1 _1213_/D sky130_fd_sc_hd__inv_2
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input222_A wr_data[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0914__A _0914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1745__A _1745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output539_A _2086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1480__A _1487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2151_ _2155_/CLK _2151_/D vssd1 vssd1 vccd1 vccd1 _2151_/Q sky130_fd_sc_hd__dfxtp_4
X_2082_ _2149_/CLK _2082_/D vssd1 vssd1 vccd1 vccd1 _2082_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1102_ _1102_/A vssd1 vssd1 vccd1 vccd1 _1102_/X sky130_fd_sc_hd__clkbuf_2
X_1033_ _1733_/A _2151_/Q _1745_/A vssd1 vssd1 vccd1 vccd1 _1034_/A sky130_fd_sc_hd__and3_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1935_ _1934_/X _0925_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1935_/X sky130_fd_sc_hd__mux2_2
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1866_ _1865_/X _1316_/Y _2013_/S vssd1 vssd1 vccd1 vccd1 _1866_/X sky130_fd_sc_hd__mux2_1
Xinput72 dout0_to_sram[27] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_6
Xinput61 dout0_to_sram[17] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_8
Xinput50 core0_data_print[7] vssd1 vssd1 vccd1 vccd1 _1089_/B sky130_fd_sc_hd__clkbuf_2
X_1797_ _1188_/Y _1796_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1797_/X sky130_fd_sc_hd__mux2_8
Xinput94 la_data_in[18] vssd1 vssd1 vccd1 vccd1 _1698_/A sky130_fd_sc_hd__buf_4
Xinput83 dout0_to_sram[8] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__buf_12
XFILLER_107_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater651 _1954_/S vssd1 vssd1 vccd1 vccd1 _2010_/S sky130_fd_sc_hd__buf_8
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1429__A2 _1422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input172_A la_data_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_134_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1365__A1 _2115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A core0_data_print[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output391_A _1717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output489_A _2041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1720_ _1720_/A vssd1 vssd1 vccd1 vccd1 _1720_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ _1767_/X _2134_/D vssd1 vssd1 vccd1 vccd1 _2134_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2065_ _1767_/X _2065_/D vssd1 vssd1 vccd1 vccd1 _2065_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2021__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1016_ _1016_/A vssd1 vssd1 vccd1 vccd1 _1016_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1918_ _1917_/X _1918_/A1 _1934_/S vssd1 vssd1 vccd1 vccd1 _1918_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1849_ _1848_/X input5/X _1942_/S vssd1 vssd1 vccd1 vccd1 _1849_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1994__S _2010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0911__B _1708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput240 wr_data[37] vssd1 vssd1 vccd1 vccd1 _1909_/A1 sky130_fd_sc_hd__buf_2
XFILLER_88_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput251 wr_data[47] vssd1 vssd1 vccd1 vccd1 _1949_/A1 sky130_fd_sc_hd__buf_2
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2044__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput262 wr_data[57] vssd1 vssd1 vccd1 vccd1 _1989_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput284 wr_data[77] vssd1 vssd1 vccd1 vccd1 _1940_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput273 wr_data[67] vssd1 vssd1 vccd1 vccd1 _1900_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput295 wr_data[87] vssd1 vssd1 vccd1 vccd1 _1980_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1510__A1 _2080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output404_A _1729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1703_ _1703_/A vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1553__660 vssd1 vssd1 vccd1 vccd1 _1553__660/HI la_data_out[1] sky130_fd_sc_hd__conb_1
XFILLER_101_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1496_ _2070_/Q _1493_/X input60/X _1494_/X vssd1 vssd1 vccd1 vccd1 _2070_/D sky130_fd_sc_hd__a22o_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2117_ _2149_/CLK _2117_/D vssd1 vssd1 vccd1 vccd1 _2117_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ _2155_/CLK _2048_/D vssd1 vssd1 vccd1 vccd1 _2048_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1099__B _1099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_129_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2067__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input135_A la_data_in[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1989__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input302_A wr_data[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_127_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1753__A _1753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1350_ _1349_/A _1339_/Y _1349_/Y _1339_/A vssd1 vssd1 vccd1 vccd1 _1350_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output521_A _2070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output619_A _1102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1281_ _1284_/A vssd1 vssd1 vccd1 vccd1 _1319_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1899__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1495__B1 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0996_ _0996_/A vssd1 vssd1 vccd1 vccd1 _0996_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput511 _2061_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[39] sky130_fd_sc_hd__buf_2
Xoutput500 _2051_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[29] sky130_fd_sc_hd__buf_2
Xoutput533 _2081_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[59] sky130_fd_sc_hd__buf_2
Xoutput522 _2071_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[49] sky130_fd_sc_hd__buf_2
XFILLER_133_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput544 _2091_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[69] sky130_fd_sc_hd__buf_2
Xoutput577 _2121_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[99] sky130_fd_sc_hd__buf_2
Xoutput566 _2111_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[89] sky130_fd_sc_hd__buf_2
Xoutput555 _2101_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[79] sky130_fd_sc_hd__buf_2
XFILLER_115_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1548_ _2110_/Q _1519_/A input69/X _1520_/A vssd1 vssd1 vccd1 vccd1 _2110_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput599 _1761_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[27] sky130_fd_sc_hd__buf_2
Xoutput588 _1751_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[17] sky130_fd_sc_hd__buf_2
X_1479_ _1486_/A vssd1 vssd1 vccd1 vccd1 _1479_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_131_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input252_A wr_data[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1477__B1 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1748__A _1748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0850_ _0875_/C vssd1 vssd1 vccd1 vccd1 _0873_/C sky130_fd_sc_hd__inv_2
XANTENNA_output471_A _2140_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output569_A _2113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1401__B1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1402_ _2137_/Q _1396_/X input63/X _1397_/X vssd1 vssd1 vccd1 vccd1 _2137_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1333_ input9/X _1320_/Y _1332_/X vssd1 vssd1 vccd1 vccd1 _1333_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1264_ input3/X _1252_/Y _1274_/B vssd1 vssd1 vccd1 vccd1 _1264_/X sky130_fd_sc_hd__o21a_1
Xinput4 addr_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
XFILLER_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1665__772 vssd1 vssd1 vccd1 vccd1 _1665__772/HI la_data_out[114] sky130_fd_sc_hd__conb_1
XFILLER_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1195_ _1195_/A _1195_/B vssd1 vssd1 vccd1 vccd1 _1206_/B sky130_fd_sc_hd__or2_1
XFILLER_25_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0979_ _1732_/A _1724_/A vssd1 vssd1 vccd1 vccd1 _0980_/A sky130_fd_sc_hd__and2_1
XFILLER_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput341 _1681_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[1] sky130_fd_sc_hd__buf_2
Xoutput330 _1680_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[0] sky130_fd_sc_hd__buf_2
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput352 _1032_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[10] sky130_fd_sc_hd__buf_2
Xoutput374 _1072_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[30] sky130_fd_sc_hd__buf_2
Xoutput396 _1721_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[21] sky130_fd_sc_hd__buf_2
XFILLER_86_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput363 _1052_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[20] sky130_fd_sc_hd__buf_2
Xoutput385 _1711_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[11] sky130_fd_sc_hd__buf_2
XFILLER_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2105__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input63_A dout0_to_sram[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1934__A1 _1934_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1162__A2 _1150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1649__756 vssd1 vssd1 vccd1 vccd1 _1649__756/HI la_data_out[97] sky130_fd_sc_hd__conb_1
XFILLER_76_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output317_A _1869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1870__A0 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1951_ _1950_/X _0942_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1951_/X sky130_fd_sc_hd__mux2_4
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0902_ _0902_/A vssd1 vssd1 vccd1 vccd1 _0902_/X sky130_fd_sc_hd__clkbuf_1
X_1882_ _1349_/A _1352_/X _1882_/S vssd1 vssd1 vccd1 vccd1 _1882_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2128__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1316_ _1319_/C _1314_/B _1315_/Y vssd1 vssd1 vccd1 vccd1 _1316_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1247_ _1263_/A vssd1 vssd1 vccd1 vccd1 _1252_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1178_ _1186_/A vssd1 vssd1 vccd1 vccd1 _1212_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input215_A wr_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1997__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1852__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0914__B _0930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0930__A _0930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output434_A _1999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1761__A _1761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2150_ _2155_/CLK _2150_/D vssd1 vssd1 vccd1 vccd1 _2150_/Q sky130_fd_sc_hd__dfxtp_1
X_2081_ _2149_/CLK _2081_/D vssd1 vssd1 vccd1 vccd1 _2081_/Q sky130_fd_sc_hd__dfxtp_2
X_1101_ _2019_/Q _1101_/B vssd1 vssd1 vccd1 vccd1 _1102_/A sky130_fd_sc_hd__and2_1
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1032_ _1032_/A vssd1 vssd1 vccd1 vccd1 _1032_/X sky130_fd_sc_hd__buf_4
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1934_ _1933_/X _1934_/A1 _1934_/S vssd1 vssd1 vccd1 vccd1 _1934_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1001__A _1001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput40 core0_data_print[27] vssd1 vssd1 vccd1 vccd1 _1129_/B sky130_fd_sc_hd__clkbuf_1
X_1865_ _1864_/X _1318_/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1865_/X sky130_fd_sc_hd__mux2_1
Xinput62 dout0_to_sram[18] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_6
Xinput73 dout0_to_sram[28] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_6
XANTENNA__0840__A _2154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1796_ _1795_/X _1684_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1796_/X sky130_fd_sc_hd__mux2_1
Xinput51 core0_data_print[8] vssd1 vssd1 vccd1 vccd1 _1091_/B sky130_fd_sc_hd__clkbuf_2
Xinput84 dout0_to_sram[9] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__buf_12
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput95 la_data_in[19] vssd1 vssd1 vccd1 vccd1 _1699_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater652 _1942_/S vssd1 vssd1 vccd1 vccd1 _1954_/S sky130_fd_sc_hd__buf_6
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1834__A0 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input165_A la_data_in[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1570__677 vssd1 vssd1 vccd1 vccd1 _1570__677/HI la_data_out[18] sky130_fd_sc_hd__conb_1
XFILLER_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0909__B _0909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input26_A core0_data_print[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1756__A _1756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output384_A _1710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output551_A _2097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2002__A0 _2001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_113_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2133_ _1767_/X _2133_/D vssd1 vssd1 vccd1 vccd1 _2133_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2064_ _1767_/X _2064_/D vssd1 vssd1 vccd1 vccd1 _2064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1015_ _1733_/A _2151_/Q _1736_/A vssd1 vssd1 vccd1 vccd1 _1016_/A sky130_fd_sc_hd__and3_1
XANTENNA__1816__A0 _1223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1917_ _1916_/X _1917_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1917_/X sky130_fd_sc_hd__mux2_2
XFILLER_135_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1848_ _1847_/X _1283_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1848_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1779_ _1156_/X _1778_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1779_/X sky130_fd_sc_hd__mux2_8
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1283__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_127_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input282_A wr_data[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput252 wr_data[48] vssd1 vssd1 vccd1 vccd1 _1953_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput241 wr_data[38] vssd1 vssd1 vccd1 vccd1 _1913_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput230 wr_data[28] vssd1 vssd1 vccd1 vccd1 _2002_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput263 wr_data[58] vssd1 vssd1 vccd1 vccd1 _1993_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput296 wr_data[88] vssd1 vssd1 vccd1 vccd1 _1984_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput285 wr_data[78] vssd1 vssd1 vccd1 vccd1 _1944_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput274 wr_data[68] vssd1 vssd1 vccd1 vccd1 _1904_/A1 sky130_fd_sc_hd__buf_2
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output599_A _1761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1702_ _1702_/A vssd1 vssd1 vccd1 vccd1 _1702_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1495_ _2069_/Q _1493_/X input59/X _1494_/X vssd1 vssd1 vccd1 vccd1 _2069_/D sky130_fd_sc_hd__a22o_1
XFILLER_4_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2116_ _2149_/CLK _2116_/D vssd1 vssd1 vccd1 vccd1 _2116_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2047_ _2155_/CLK _2047_/D vssd1 vssd1 vccd1 vccd1 _2047_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input128_A la_data_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0922__B _0930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input93_A la_data_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1576__683 vssd1 vssd1 vccd1 vccd1 _1576__683/HI la_data_out[24] sky130_fd_sc_hd__conb_1
XFILLER_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output347_A _1687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1280_ input5/X vssd1 vssd1 vccd1 vccd1 _1284_/A sky130_fd_sc_hd__inv_2
XFILLER_95_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output514_A _2063_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1495__A1 _2069_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0995_ _1732_/A _1728_/A vssd1 vssd1 vccd1 vccd1 _0996_/A sky130_fd_sc_hd__and2_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_117_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput501 _2024_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[2] sky130_fd_sc_hd__buf_2
Xoutput534 _2027_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[5] sky130_fd_sc_hd__buf_2
Xoutput545 _2028_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[6] sky130_fd_sc_hd__buf_2
Xoutput523 _2026_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[4] sky130_fd_sc_hd__buf_2
Xoutput512 _2025_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput556 _2029_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[7] sky130_fd_sc_hd__buf_2
Xoutput567 _2030_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[8] sky130_fd_sc_hd__buf_2
Xoutput578 _2031_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_99_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1547_ _2109_/Q _1519_/A input68/X _1520_/A vssd1 vssd1 vccd1 vccd1 _2109_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput589 _1752_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[18] sky130_fd_sc_hd__buf_2
XFILLER_115_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1478_ _2058_/Q _1470_/X input79/X _1473_/X vssd1 vssd1 vccd1 vccd1 _2058_/D sky130_fd_sc_hd__a22o_1
XFILLER_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1238__A1 _1235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2034__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1610__717 vssd1 vssd1 vccd1 vccd1 _1610__717/HI la_data_out[58] sky130_fd_sc_hd__conb_1
XFILLER_2_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input245_A wr_data[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1477__B2 _1473_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1229__A1 _1223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1401__A1 _2136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1401__B2 _1397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output464_A _2133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1764__A _1764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1401_ _2136_/Q _1396_/X input62/X _1397_/X vssd1 vssd1 vccd1 vccd1 _2136_/D sky130_fd_sc_hd__a22o_1
XANTENNA_output631_A _1124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1332_ _1343_/A _1343_/C vssd1 vssd1 vccd1 vccd1 _1332_/X sky130_fd_sc_hd__or2_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1263_ _1263_/A _1265_/A _1263_/C vssd1 vssd1 vccd1 vccd1 _1274_/B sky130_fd_sc_hd__or3_1
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput5 addr_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
XFILLER_64_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1194_ _1195_/A _1193_/B _1204_/B vssd1 vssd1 vccd1 vccd1 _1194_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2057__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0978_ _0978_/A vssd1 vssd1 vccd1 vccd1 _0978_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput342 _1682_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[2] sky130_fd_sc_hd__buf_2
XFILLER_133_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput331 _1690_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[10] sky130_fd_sc_hd__buf_2
Xoutput353 _1034_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[11] sky130_fd_sc_hd__buf_2
Xoutput320 _1887_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[19] sky130_fd_sc_hd__buf_2
XFILLER_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput375 _1074_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[31] sky130_fd_sc_hd__buf_2
Xoutput364 _1054_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[21] sky130_fd_sc_hd__buf_2
Xoutput386 _1712_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[12] sky130_fd_sc_hd__buf_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput397 _1722_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[22] sky130_fd_sc_hd__buf_2
XFILLER_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input195_A wr_data[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1395__B1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input56_A dout0_to_sram[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0928__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1759__A _1759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1950_ _1949_/X _1950_/A1 _2010_/S vssd1 vssd1 vccd1 vccd1 _1950_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0901_ _0901_/A _0909_/B vssd1 vssd1 vccd1 vccd1 _0902_/A sky130_fd_sc_hd__and2_2
X_1881_ _1348_/Y _1880_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__mux2_4
XFILLER_115_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1386__B1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1315_ _1327_/B vssd1 vssd1 vccd1 vccd1 _1315_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1246_ input2/X vssd1 vssd1 vccd1 vccd1 _1263_/A sky130_fd_sc_hd__inv_2
XFILLER_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1177_ _1177_/A vssd1 vssd1 vccd1 vccd1 _1186_/A sky130_fd_sc_hd__inv_2
XFILLER_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1861__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1377__B1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input110_A la_data_in[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input208_A wr_data[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1616__723 vssd1 vssd1 vccd1 vccd1 _1616__723/HI la_data_out[64] sky130_fd_sc_hd__conb_1
XFILLER_125_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1368__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0930__B _0930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output427_A _1971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1100_ _1100_/A vssd1 vssd1 vccd1 vccd1 _1100_/X sky130_fd_sc_hd__buf_2
XFILLER_93_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2080_ _1767_/X _2080_/D vssd1 vssd1 vccd1 vccd1 _2080_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1031_ _1733_/A _2151_/Q _1744_/A vssd1 vssd1 vccd1 vccd1 _1032_/A sky130_fd_sc_hd__and3_1
XFILLER_62_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1843__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1933_ _1932_/X _1933_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1933_/X sky130_fd_sc_hd__mux2_4
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1001__B _1009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 core0_data_print[18] vssd1 vssd1 vccd1 vccd1 _1111_/B sky130_fd_sc_hd__clkbuf_2
X_1864_ input8/X _1321_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1864_/X sky130_fd_sc_hd__mux2_1
Xinput41 core0_data_print[28] vssd1 vssd1 vccd1 vccd1 _1131_/B sky130_fd_sc_hd__buf_2
Xinput63 dout0_to_sram[19] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_6
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput52 core0_data_print[9] vssd1 vssd1 vccd1 vccd1 _1093_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__0840__B _2152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1795_ _1794_/X _1177_/A _1922_/S vssd1 vssd1 vccd1 vccd1 _1795_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput74 dout0_to_sram[29] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_6
Xinput96 la_data_in[1] vssd1 vssd1 vccd1 vccd1 _1681_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 la_data_in[0] vssd1 vssd1 vccd1 vccd1 _1680_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1531__B1 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater653 _1938_/S vssd1 vssd1 vccd1 vccd1 _1942_/S sky130_fd_sc_hd__buf_6
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1229_ _1223_/A _1216_/Y _1239_/B vssd1 vssd1 vccd1 vccd1 _1229_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_119_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input158_A la_data_in[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1522__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input19_A addr_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1801__S _1922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1825__A1 _1235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_129_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2118__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0941__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output377_A _1020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2002__A1 _2002_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output544_A _2091_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1513__B1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _2149_/CLK _2132_/D vssd1 vssd1 vccd1 vccd1 _2132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2063_ _2155_/CLK _2063_/D vssd1 vssd1 vccd1 vccd1 _2063_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1014_ _1014_/A vssd1 vssd1 vccd1 vccd1 _1014_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1916_ _0910_/X _1916_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1916_/X sky130_fd_sc_hd__mux2_4
XFILLER_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1847_ _1846_/X _1286_/Y _2012_/S vssd1 vssd1 vccd1 vccd1 _1847_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1778_ _1777_/X _1681_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1778_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1504__B1 input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input275_A wr_data[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput220 wr_data[19] vssd1 vssd1 vccd1 vccd1 _1966_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput231 wr_data[29] vssd1 vssd1 vccd1 vccd1 _2006_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput253 wr_data[49] vssd1 vssd1 vccd1 vccd1 _1957_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput242 wr_data[39] vssd1 vssd1 vccd1 vccd1 _1917_/A1 sky130_fd_sc_hd__buf_2
Xinput286 wr_data[79] vssd1 vssd1 vccd1 vccd1 _1948_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput264 wr_data[59] vssd1 vssd1 vccd1 vccd1 _1997_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput297 wr_data[89] vssd1 vssd1 vccd1 vccd1 _1988_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_76_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput275 wr_data[69] vssd1 vssd1 vccd1 vccd1 _1908_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output494_A _2045_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__2090__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1701_ _1701_/A vssd1 vssd1 vccd1 vccd1 _1701_/X sky130_fd_sc_hd__buf_2
XANTENNA__1982__A0 _1981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1494_ _1508_/A vssd1 vssd1 vccd1 vccd1 _1494_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1007__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2115_ _1767_/X _2115_/D vssd1 vssd1 vccd1 vccd1 _2115_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2046_ _2149_/CLK _2046_/D vssd1 vssd1 vccd1 vccd1 _2046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input86_A la_data_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_122_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater657_A _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0994_ _0994_/A vssd1 vssd1 vccd1 vccd1 _0994_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput502 _2052_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[30] sky130_fd_sc_hd__buf_2
Xoutput513 _2062_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[40] sky130_fd_sc_hd__buf_2
XFILLER_132_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput535 _2082_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[60] sky130_fd_sc_hd__buf_2
Xoutput524 _2072_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[50] sky130_fd_sc_hd__buf_2
Xoutput546 _2092_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[70] sky130_fd_sc_hd__buf_2
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1546_ _2108_/Q _1540_/X input67/X _1541_/X vssd1 vssd1 vccd1 vccd1 _2108_/D sky130_fd_sc_hd__a22o_1
Xoutput557 _2102_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[80] sky130_fd_sc_hd__buf_2
XFILLER_5_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput568 _2112_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[90] sky130_fd_sc_hd__buf_2
XFILLER_115_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput579 _1733_/X vssd1 vssd1 vccd1 vccd1 read_enable_to_Elpis sky130_fd_sc_hd__buf_2
XFILLER_99_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1477_ _2057_/Q _1470_/X input78/X _1473_/X vssd1 vssd1 vccd1 vccd1 _2057_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2029_ _2155_/CLK _2029_/D vssd1 vssd1 vccd1 vccd1 _2029_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_24_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1946__A0 _1945_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input238_A wr_data[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input140_A la_data_in[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1477__A2 _1470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1401__A2 _1396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1400_ _2135_/Q _1396_/X input61/X _1397_/X vssd1 vssd1 vccd1 vccd1 _2135_/D sky130_fd_sc_hd__a22o_1
XANTENNA_output457_A _2127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output624_A _1112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1331_ _1343_/A _1329_/B _1330_/Y vssd1 vssd1 vccd1 vccd1 _1331_/Y sky130_fd_sc_hd__a21oi_1
X_1262_ _1265_/A _1260_/B _1261_/Y vssd1 vssd1 vccd1 vccd1 _1262_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput6 addr_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_4
XFILLER_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1193_ _1212_/B _1193_/B vssd1 vssd1 vccd1 vccd1 _1204_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0977_ _0977_/A _0993_/B vssd1 vssd1 vccd1 vccd1 _0978_/A sky130_fd_sc_hd__and2_1
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput310 _1773_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[0] sky130_fd_sc_hd__buf_2
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput343 _1683_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[3] sky130_fd_sc_hd__buf_2
XFILLER_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput321 _1779_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[1] sky130_fd_sc_hd__buf_2
Xoutput332 _1691_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[11] sky130_fd_sc_hd__buf_2
Xoutput365 _1056_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[22] sky130_fd_sc_hd__buf_2
Xoutput354 _1036_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[12] sky130_fd_sc_hd__buf_2
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput376 _1018_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[3] sky130_fd_sc_hd__buf_2
Xoutput387 _1713_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[13] sky130_fd_sc_hd__buf_2
Xoutput398 _1723_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[23] sky130_fd_sc_hd__buf_2
X_1529_ _2095_/Q _1526_/X input84/X _1527_/X vssd1 vssd1 vccd1 vccd1 _2095_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2151__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input188_A wr_data[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input49_A core0_data_print[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1804__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0928__B _1712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1105__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0900_ _0900_/A vssd1 vssd1 vccd1 vccd1 _0900_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1880_ _1879_/X _1698_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1880_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output574_A _2118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1386__A1 _2125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1314_ _1322_/A _1314_/B vssd1 vssd1 vccd1 vccd1 _1327_/B sky130_fd_sc_hd__or2_1
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1015__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1245_ _1235_/A _1233_/Y _1254_/B vssd1 vssd1 vccd1 vccd1 _1245_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2024__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1176_ _1168_/B _1165_/Y _1186_/B vssd1 vssd1 vccd1 vccd1 _1176_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0854__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1685__A _1685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1377__A1 _2118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input103_A la_data_in[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1655__762 vssd1 vssd1 vccd1 vccd1 _1655__762/HI la_data_out[104] sky130_fd_sc_hd__conb_1
XANTENNA__1368__A1 _2116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2047__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1030_ _1030_/A vssd1 vssd1 vccd1 vccd1 _1030_/X sky130_fd_sc_hd__buf_2
XFILLER_62_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1932_ _0927_/X _1932_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1932_/X sky130_fd_sc_hd__mux2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1863_ _1311_/X _1862_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1863_/X sky130_fd_sc_hd__mux2_4
Xinput31 core0_data_print[19] vssd1 vssd1 vccd1 vccd1 _1113_/B sky130_fd_sc_hd__clkbuf_4
Xinput20 addr_in[9] vssd1 vssd1 vccd1 vccd1 _1235_/A sky130_fd_sc_hd__buf_4
Xinput53 dout0_to_sram[0] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_12
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput64 dout0_to_sram[1] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_8
Xinput42 core0_data_print[29] vssd1 vssd1 vccd1 vccd1 _1133_/B sky130_fd_sc_hd__buf_2
X_1794_ _1793_/X _1181_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1794_/X sky130_fd_sc_hd__mux2_1
Xinput75 dout0_to_sram[2] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_12
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput97 la_data_in[2] vssd1 vssd1 vccd1 vccd1 _1682_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput86 la_data_in[10] vssd1 vssd1 vccd1 vccd1 _1690_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0849__A _2152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1531__A1 _2097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater654 _1958_/S vssd1 vssd1 vccd1 vccd1 _1938_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_72_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1228_ _1228_/A _1228_/B vssd1 vssd1 vccd1 vccd1 _1239_/B sky130_fd_sc_hd__or2_1
XFILLER_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1159_ _1168_/A vssd1 vssd1 vccd1 vccd1 _1175_/A sky130_fd_sc_hd__inv_2
X_1598__705 vssd1 vssd1 vccd1 vccd1 _1598__705/HI la_data_out[46] sky130_fd_sc_hd__conb_1
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1639__746 vssd1 vssd1 vccd1 vccd1 _1639__746/HI la_data_out[87] sky130_fd_sc_hd__conb_1
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1522__A1 _2090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input220_A wr_data[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0941__B _1715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_138_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output537_A _2084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1513__A1 _2083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2131_ _2149_/CLK _2131_/D vssd1 vssd1 vccd1 vccd1 _2131_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2062_ _2155_/CLK _2062_/D vssd1 vssd1 vccd1 vccd1 _2062_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1013_ _1733_/A _2151_/Q _1735_/A vssd1 vssd1 vccd1 vccd1 _1014_/A sky130_fd_sc_hd__and3_1
XFILLER_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1915_ _1914_/X _0904_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1915_/X sky130_fd_sc_hd__mux2_4
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1846_ input5/X _1288_/X _1882_/S vssd1 vssd1 vccd1 vccd1 _1846_/X sky130_fd_sc_hd__mux2_1
X_1777_ _1776_/X _1150_/A _1922_/S vssd1 vssd1 vccd1 vccd1 _1777_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1504__A1 _2076_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1902__S _1958_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1440__B1 _2032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input170_A la_data_in[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input268_A wr_data[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput210 wr_data[125] vssd1 vssd1 vccd1 vccd1 _1001_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input31_A core0_data_print[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput221 wr_data[1] vssd1 vssd1 vccd1 vccd1 _1894_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput232 wr_data[2] vssd1 vssd1 vccd1 vccd1 _1898_/A1 sky130_fd_sc_hd__buf_4
Xinput243 wr_data[3] vssd1 vssd1 vccd1 vccd1 _1902_/A1 sky130_fd_sc_hd__buf_2
Xinput254 wr_data[4] vssd1 vssd1 vccd1 vccd1 _1906_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput287 wr_data[7] vssd1 vssd1 vccd1 vccd1 _1918_/A1 sky130_fd_sc_hd__buf_2
XFILLER_84_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput276 wr_data[6] vssd1 vssd1 vccd1 vccd1 _1914_/A1 sky130_fd_sc_hd__buf_2
Xinput265 wr_data[5] vssd1 vssd1 vccd1 vccd1 _1910_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__1812__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput298 wr_data[8] vssd1 vssd1 vccd1 vccd1 _1922_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1113__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output487_A _2039_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1700_ _1700_/A vssd1 vssd1 vccd1 vccd1 _1700_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1982__A1 _1982_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1493_ _1507_/A vssd1 vssd1 vccd1 vccd1 _1493_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1007__B _1731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1498__B1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2114_ _1767_/X _2114_/D vssd1 vssd1 vccd1 vccd1 _2114_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1023__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2045_ _2155_/CLK _2045_/D vssd1 vssd1 vccd1 vccd1 _2045_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1560__667 vssd1 vssd1 vccd1 vccd1 _1560__667/HI la_data_out[8] sky130_fd_sc_hd__conb_1
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1829_ _1828_/X _1251_/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1829_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1693__A _1693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2108__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1489__B1 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_85_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_13_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_110_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1413__B1 input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1964__A1 _1964_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input79_A dout0_to_sram[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1807__S _1922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output402_A _1727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0993_ _0993_/A _0993_/B vssd1 vssd1 vccd1 vccd1 _0994_/A sky130_fd_sc_hd__and2_1
XFILLER_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput536 _2083_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[61] sky130_fd_sc_hd__buf_2
Xoutput525 _2073_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[51] sky130_fd_sc_hd__buf_2
Xoutput503 _2053_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[31] sky130_fd_sc_hd__buf_2
Xoutput514 _2063_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[41] sky130_fd_sc_hd__buf_2
XFILLER_132_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput569 _2113_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[91] sky130_fd_sc_hd__buf_2
X_1545_ _2107_/Q _1540_/X input66/X _1541_/X vssd1 vssd1 vccd1 vccd1 _2107_/D sky130_fd_sc_hd__a22o_1
Xoutput558 _2103_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[81] sky130_fd_sc_hd__buf_2
XFILLER_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput547 _2093_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[71] sky130_fd_sc_hd__buf_2
XFILLER_115_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1476_ _2056_/Q _1470_/X input75/X _1473_/X vssd1 vssd1 vccd1 vccd1 _2056_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2028_ _2155_/CLK _2028_/D vssd1 vssd1 vccd1 vccd1 _2028_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1688__A _1688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1946__A1 _1946_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input133_A la_data_in[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2080__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1882__A0 _1349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input300_A wr_data[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_5_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output352_A _1032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1330_ _1341_/B vssd1 vssd1 vccd1 vccd1 _1330_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1261_ _1272_/B vssd1 vssd1 vccd1 vccd1 _1261_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1192_ _1195_/A _1191_/B _1202_/B vssd1 vssd1 vccd1 vccd1 _1192_/Y sky130_fd_sc_hd__a21boi_1
Xinput7 addr_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
XFILLER_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1301__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0976_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0993_/B sky130_fd_sc_hd__buf_2
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_133_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput333 _1692_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[12] sky130_fd_sc_hd__buf_2
X_1672__779 vssd1 vssd1 vccd1 vccd1 _1672__779/HI la_data_out[121] sky130_fd_sc_hd__conb_1
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput322 _1785_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[2] sky130_fd_sc_hd__buf_2
Xoutput344 _1684_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[4] sky130_fd_sc_hd__buf_2
Xoutput311 _1833_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[10] sky130_fd_sc_hd__buf_2
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput366 _1058_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[23] sky130_fd_sc_hd__buf_2
Xoutput377 _1020_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[4] sky130_fd_sc_hd__buf_2
Xoutput355 _1038_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[13] sky130_fd_sc_hd__buf_2
Xoutput399 _1724_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[24] sky130_fd_sc_hd__buf_2
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1528_ _2094_/Q _1526_/X input83/X _1527_/X vssd1 vssd1 vccd1 vccd1 _2094_/D sky130_fd_sc_hd__a22o_1
Xoutput388 _1714_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[14] sky130_fd_sc_hd__buf_2
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1459_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1864__A0 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1566__673 vssd1 vssd1 vccd1 vccd1 _1566__673/HI la_data_out[14] sky130_fd_sc_hd__conb_1
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1910__S _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input250_A wr_data[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1105__B _1105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1820__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1121__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0960__A _0960_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1313_ _1322_/A vssd1 vssd1 vccd1 vccd1 _1319_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1244_ _1244_/A _1244_/B vssd1 vssd1 vccd1 vccd1 _1254_/B sky130_fd_sc_hd__or2_1
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1015__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1846__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1175_ _1175_/A _1175_/B _1175_/C vssd1 vssd1 vccd1 vccd1 _1186_/B sky130_fd_sc_hd__or3_1
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1031__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1600__707 vssd1 vssd1 vccd1 vccd1 _1600__707/HI la_data_out[48] sky130_fd_sc_hd__conb_1
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0959_ _0959_/A vssd1 vssd1 vccd1 vccd1 _0959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1905__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input298_A wr_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2014__A0 _2013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input61_A dout0_to_sram[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1815__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0939__B _0951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1828__A0 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1931_ _1930_/X _0921_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1931_/X sky130_fd_sc_hd__mux2_1
X_1862_ _1861_/X _1695_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1862_/X sky130_fd_sc_hd__mux2_1
Xinput21 core0_data_print[0] vssd1 vssd1 vccd1 vccd1 _1075_/B sky130_fd_sc_hd__buf_4
XANTENNA__2005__A0 _2004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput10 addr_in[18] vssd1 vssd1 vccd1 vccd1 _1336_/A sky130_fd_sc_hd__buf_2
XFILLER_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput54 dout0_to_sram[10] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_16
Xinput32 core0_data_print[1] vssd1 vssd1 vccd1 vccd1 _1077_/B sky130_fd_sc_hd__buf_2
Xinput43 core0_data_print[2] vssd1 vssd1 vccd1 vccd1 _1079_/B sky130_fd_sc_hd__clkbuf_1
X_1793_ _1792_/X _1183_/Y _2012_/S vssd1 vssd1 vccd1 vccd1 _1793_/X sky130_fd_sc_hd__mux2_1
Xinput87 la_data_in[11] vssd1 vssd1 vccd1 vccd1 _1691_/A sky130_fd_sc_hd__buf_4
XFILLER_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput76 dout0_to_sram[30] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_6
Xinput65 dout0_to_sram[20] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_6
Xinput98 la_data_in[32] vssd1 vssd1 vccd1 vccd1 _1700_/A sky130_fd_sc_hd__buf_6
XFILLER_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2141__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater655 _1958_/S vssd1 vssd1 vccd1 vccd1 _1922_/S sky130_fd_sc_hd__buf_6
X_1227_ _1232_/A _1225_/B _1226_/Y vssd1 vssd1 vccd1 vccd1 _1227_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1158_ _1168_/A _1168_/C _1157_/Y vssd1 vssd1 vccd1 vccd1 _1158_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1089_ _2019_/Q _1089_/B vssd1 vssd1 vccd1 vccd1 _1090_/A sky130_fd_sc_hd__and2_1
XFILLER_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1696__A _1696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1678__785 vssd1 vssd1 vccd1 vccd1 _1678__785/HI la_data_out[127] sky130_fd_sc_hd__conb_1
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input213_A wr_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_112_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output432_A _1991_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2130_ _2149_/CLK _2130_/D vssd1 vssd1 vccd1 vccd1 _2130_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2061_ _2155_/CLK _2061_/D vssd1 vssd1 vccd1 vccd1 _2061_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1012_ _1012_/A vssd1 vssd1 vccd1 vccd1 _1012_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1914_ _1913_/X _1914_/A1 _1934_/S vssd1 vssd1 vccd1 vccd1 _1914_/X sky130_fd_sc_hd__mux2_1
X_1845_ _1279_/Y _1844_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1845_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1776_ _1775_/X _1154_/A _2013_/S vssd1 vssd1 vccd1 vccd1 _1776_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1606__713 vssd1 vssd1 vccd1 vccd1 _1606__713/HI la_data_out[54] sky130_fd_sc_hd__conb_1
XFILLER_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2037__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1440__A1 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input163_A la_data_in[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput211 wr_data[126] vssd1 vssd1 vccd1 vccd1 _1005_/A sky130_fd_sc_hd__buf_4
Xinput200 wr_data[116] vssd1 vssd1 vccd1 vccd1 _0964_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput222 wr_data[20] vssd1 vssd1 vccd1 vccd1 _1970_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput244 wr_data[40] vssd1 vssd1 vccd1 vccd1 _1921_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xinput233 wr_data[30] vssd1 vssd1 vccd1 vccd1 _2010_/A1 sky130_fd_sc_hd__buf_2
Xinput277 wr_data[70] vssd1 vssd1 vccd1 vccd1 _1912_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput266 wr_data[60] vssd1 vssd1 vccd1 vccd1 _2001_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput288 wr_data[80] vssd1 vssd1 vccd1 vccd1 _1952_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput255 wr_data[50] vssd1 vssd1 vccd1 vccd1 _1961_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input24_A core0_data_print[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput299 wr_data[90] vssd1 vssd1 vccd1 vccd1 _1992_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1259__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1113__B _1113_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output382_A _1030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output647_A _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1492_ _2068_/Q _1486_/X input58/X _1487_/X vssd1 vssd1 vccd1 vccd1 _2068_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1498__A1 _2072_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2113_ _1767_/X _2113_/D vssd1 vssd1 vccd1 vccd1 _2113_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2044_ _2155_/CLK _2044_/D vssd1 vssd1 vccd1 vccd1 _2044_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1023__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1828_ input2/X _1253_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1828_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1759_ _1759_/A vssd1 vssd1 vccd1 vccd1 _1759_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_89_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1913__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2020__D _2154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1413__A1 _2144_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input280_A wr_data[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1823__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0947__B _0951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output597_A _1759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0992_ _0992_/A vssd1 vssd1 vccd1 vccd1 _0992_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput526 _2074_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[52] sky130_fd_sc_hd__buf_2
Xoutput515 _2064_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[42] sky130_fd_sc_hd__buf_2
Xoutput504 _2054_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[32] sky130_fd_sc_hd__buf_2
Xoutput537 _2084_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[62] sky130_fd_sc_hd__buf_2
Xoutput559 _2104_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[82] sky130_fd_sc_hd__buf_2
Xoutput548 _2094_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[72] sky130_fd_sc_hd__buf_2
X_1544_ _2106_/Q _1540_/X input65/X _1541_/X vssd1 vssd1 vccd1 vccd1 _2106_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_113_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1475_ _2055_/Q _1470_/X input64/X _1473_/X vssd1 vssd1 vccd1 vccd1 _2055_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2027_ _2155_/CLK _2027_/D vssd1 vssd1 vccd1 vccd1 _2027_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1908__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input126_A la_data_in[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input91_A la_data_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1398__B1 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1818__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1119__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0958__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1260_ _1265_/A _1260_/B vssd1 vssd1 vccd1 vccd1 _1272_/B sky130_fd_sc_hd__or2_1
XFILLER_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1191_ _1195_/A _1191_/B vssd1 vssd1 vccd1 vccd1 _1202_/B sky130_fd_sc_hd__or2_1
Xinput8 addr_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_92_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1873__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0975_ _0975_/A vssd1 vssd1 vccd1 vccd1 _0975_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput312 _1839_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[11] sky130_fd_sc_hd__buf_2
XFILLER_133_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput323 _1791_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[3] sky130_fd_sc_hd__buf_2
XANTENNA__1029__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput334 _1693_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[13] sky130_fd_sc_hd__buf_2
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput367 _1060_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[24] sky130_fd_sc_hd__buf_2
Xoutput378 _1022_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[5] sky130_fd_sc_hd__buf_2
Xoutput345 _1685_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[5] sky130_fd_sc_hd__buf_2
Xoutput356 _1040_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[14] sky130_fd_sc_hd__buf_2
Xoutput389 _1715_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[15] sky130_fd_sc_hd__buf_2
X_1527_ _1541_/A vssd1 vssd1 vccd1 vccd1 _1527_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1458_ input69/X _1452_/X _2046_/Q _1453_/X vssd1 vssd1 vccd1 vccd1 _2046_/D sky130_fd_sc_hd__o22a_1
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1389_ _1389_/A vssd1 vssd1 vccd1 vccd1 _1389_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1699__A _1699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input243_A wr_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1855__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1121__B _1121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0960__B _0972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output462_A _2032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1543__B1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1312_ input8/X vssd1 vssd1 vccd1 vccd1 _1322_/A sky130_fd_sc_hd__inv_2
XFILLER_111_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1589__696 vssd1 vssd1 vccd1 vccd1 _1589__696/HI la_data_out[37] sky130_fd_sc_hd__conb_1
X_1243_ _1244_/A _1242_/B _1263_/C vssd1 vssd1 vccd1 vccd1 _1243_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_49_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1015__C _1736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1174_ _1168_/B _1162_/X _1184_/B vssd1 vssd1 vccd1 vccd1 _1174_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1312__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1031__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2070__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0958_ _1732_/A _1719_/A vssd1 vssd1 vccd1 vccd1 _0959_/A sky130_fd_sc_hd__and2_1
XFILLER_134_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0889_ _1732_/A _1703_/A vssd1 vssd1 vccd1 vccd1 _0890_/A sky130_fd_sc_hd__and2_1
XFILLER_133_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1921__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1837__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input193_A wr_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input54_A dout0_to_sram[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1525__B1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1831__S _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2093__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ _1929_/X _1930_/A1 _1938_/S vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1861_ _1860_/X input7/X _1954_/S vssd1 vssd1 vccd1 vccd1 _1861_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2005__A1 _2005_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 addr_in[19] vssd1 vssd1 vccd1 vccd1 _1349_/A sky130_fd_sc_hd__clkbuf_4
Xinput22 core0_data_print[10] vssd1 vssd1 vccd1 vccd1 _1095_/B sky130_fd_sc_hd__clkbuf_1
Xinput55 dout0_to_sram[11] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_16
XFILLER_128_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput44 core0_data_print[30] vssd1 vssd1 vccd1 vccd1 _1135_/B sky130_fd_sc_hd__buf_2
Xinput33 core0_data_print[20] vssd1 vssd1 vccd1 vccd1 _1115_/B sky130_fd_sc_hd__clkbuf_2
X_1792_ _1177_/A _1185_/X _1882_/S vssd1 vssd1 vccd1 vccd1 _1792_/X sky130_fd_sc_hd__mux2_1
Xinput77 dout0_to_sram[31] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__buf_6
Xinput66 dout0_to_sram[21] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_8
Xinput88 la_data_in[12] vssd1 vssd1 vccd1 vccd1 _1692_/A sky130_fd_sc_hd__buf_4
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput99 la_data_in[33] vssd1 vssd1 vccd1 vccd1 _1701_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1516__B1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater656 _2149_/CLK vssd1 vssd1 vccd1 vccd1 _2155_/CLK sky130_fd_sc_hd__buf_12
X_1226_ _1237_/B vssd1 vssd1 vccd1 vccd1 _1226_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1819__A1 _1223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1157_ _1168_/A _1168_/C vssd1 vssd1 vccd1 vccd1 _1157_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1088_ _1088_/A vssd1 vssd1 vccd1 vccd1 _1088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0881__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1916__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input206_A wr_data[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1994__A0 _1993_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1826__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1127__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0966__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output425_A _1967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2060_ _2155_/CLK _2060_/D vssd1 vssd1 vccd1 vccd1 _2060_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1011_ _1733_/A _2151_/Q _1734_/A vssd1 vssd1 vccd1 vccd1 _1012_/A sky130_fd_sc_hd__and3_1
XFILLER_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1913_ _1912_/X _1913_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1913_/X sky130_fd_sc_hd__mux2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1844_ _1843_/X _1692_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1844_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1775_ _1774_/X _1160_/A _2012_/S vssd1 vssd1 vccd1 vccd1 _1775_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1037__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0876__A _0876_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1209_ _1208_/A _1221_/C _1208_/Y vssd1 vssd1 vccd1 vccd1 _1209_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1645__752 vssd1 vssd1 vccd1 vccd1 _1645__752/HI la_data_out[93] sky130_fd_sc_hd__conb_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input156_A la_data_in[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput201 wr_data[117] vssd1 vssd1 vccd1 vccd1 _0968_/A sky130_fd_sc_hd__buf_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput234 wr_data[31] vssd1 vssd1 vccd1 vccd1 _2014_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput223 wr_data[21] vssd1 vssd1 vccd1 vccd1 _1974_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput212 wr_data[127] vssd1 vssd1 vccd1 vccd1 _1009_/A sky130_fd_sc_hd__buf_4
Xinput245 wr_data[41] vssd1 vssd1 vccd1 vccd1 _1925_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput278 wr_data[71] vssd1 vssd1 vccd1 vccd1 _1916_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput267 wr_data[61] vssd1 vssd1 vccd1 vccd1 _2005_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput256 wr_data[51] vssd1 vssd1 vccd1 vccd1 _1965_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput289 wr_data[81] vssd1 vssd1 vccd1 vccd1 _1956_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input17_A addr_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1967__A0 _1966_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2131__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output375_A _1074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output542_A _2089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1491_ _2067_/Q _1486_/X input57/X _1487_/X vssd1 vssd1 vccd1 vccd1 _2067_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1629__736 vssd1 vssd1 vccd1 vccd1 _1629__736/HI la_data_out[77] sky130_fd_sc_hd__conb_1
XFILLER_94_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2112_ _1767_/X _2112_/D vssd1 vssd1 vccd1 vccd1 _2112_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2043_ _2149_/CLK _2043_/D vssd1 vssd1 vccd1 vccd1 _2043_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1023__C _1740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0862__C _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1958__A0 _1957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1827_ _1245_/X _1826_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1827_/X sky130_fd_sc_hd__mux2_4
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1758_ _1758_/A vssd1 vssd1 vccd1 vccd1 _1758_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1689_ _1689_/A vssd1 vssd1 vccd1 vccd1 _1689_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input9_A addr_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1949__A0 _1948_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__2154__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input273_A wr_data[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2000__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output492_A _2043_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0991_ _1732_/A _1727_/A vssd1 vssd1 vccd1 vccd1 _0992_/A sky130_fd_sc_hd__and2_1
XFILLER_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput516 _2065_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[43] sky130_fd_sc_hd__buf_2
Xoutput505 _2055_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[33] sky130_fd_sc_hd__buf_2
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput527 _2075_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[53] sky130_fd_sc_hd__buf_2
Xoutput538 _2085_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[63] sky130_fd_sc_hd__buf_2
XFILLER_113_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1543_ _2105_/Q _1540_/X input63/X _1541_/X vssd1 vssd1 vccd1 vccd1 _2105_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput549 _2095_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[73] sky130_fd_sc_hd__buf_2
X_1474_ _2054_/Q _1470_/X input53/X _1473_/X vssd1 vssd1 vccd1 vccd1 _2054_/D sky130_fd_sc_hd__a22o_1
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2027__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0873__B _2152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2026_ _2155_/CLK _2026_/D vssd1 vssd1 vccd1 vccd1 _2026_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1924__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A la_data_in[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input84_A dout0_to_sram[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1398__B2 _1397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1398__A1 _2133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1119__B _1119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1834__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0958__B _1719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1135__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output338_A _1697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1190_ _1212_/B vssd1 vssd1 vccd1 vccd1 _1195_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output505_A _2055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0974__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 addr_in[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_18_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater655_A _1958_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0974_ _1732_/A _1723_/A vssd1 vssd1 vccd1 vccd1 _0975_/A sky130_fd_sc_hd__and2_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput324 _1797_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[4] sky130_fd_sc_hd__buf_2
XANTENNA__1029__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput335 _1694_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[14] sky130_fd_sc_hd__buf_2
Xoutput313 _1845_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[12] sky130_fd_sc_hd__buf_2
X_1526_ _1540_/A vssd1 vssd1 vccd1 vccd1 _1526_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput368 _1062_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[25] sky130_fd_sc_hd__buf_2
Xoutput346 _1686_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[6] sky130_fd_sc_hd__buf_2
Xoutput357 _1042_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[15] sky130_fd_sc_hd__buf_2
XFILLER_102_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput379 _1024_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[6] sky130_fd_sc_hd__buf_2
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1457_ input68/X _1452_/X _2045_/Q _1453_/X vssd1 vssd1 vccd1 vccd1 _2045_/D sky130_fd_sc_hd__o22a_1
XANTENNA__1045__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1388_ _2127_/Q _1382_/X input84/X _1383_/X vssd1 vssd1 vccd1 vccd1 _2127_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2009_ _2008_/X _2009_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__mux2_2
XFILLER_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1919__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_136_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_105_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input236_A wr_data[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1304__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1829__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output455_A _2125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1543__A1 _2105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output622_A _1108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1311_ input7/X _1299_/Y _1322_/B vssd1 vssd1 vccd1 vccd1 _1311_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1242_ _1244_/A _1242_/B vssd1 vssd1 vccd1 vccd1 _1263_/C sky130_fd_sc_hd__or2_1
XFILLER_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1173_ _1173_/A vssd1 vssd1 vccd1 vccd1 _1184_/B sky130_fd_sc_hd__inv_2
XFILLER_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1031__C _1744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0957_ _0957_/A vssd1 vssd1 vccd1 vccd1 _0957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0888_ _0888_/A vssd1 vssd1 vccd1 vccd1 _0888_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0879__A _0879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1509_ _2079_/Q _1507_/X input70/X _1508_/X vssd1 vssd1 vccd1 vccd1 _2079_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_109_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input186_A wr_data[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1525__A1 _2093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_79_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input47_A core0_data_print[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1662__769 vssd1 vssd1 vccd1 vccd1 _1662__769/HI la_data_out[111] sky130_fd_sc_hd__conb_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1461__B1 _2047_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1860_ _1859_/X _1304_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1860_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output572_A _2116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1791_ _1176_/X _1790_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1791_/X sky130_fd_sc_hd__mux2_1
Xinput12 addr_in[1] vssd1 vssd1 vccd1 vccd1 _1150_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput34 core0_data_print[21] vssd1 vssd1 vccd1 vccd1 _1117_/B sky130_fd_sc_hd__buf_2
Xinput23 core0_data_print[11] vssd1 vssd1 vccd1 vccd1 _1097_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_128_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput45 core0_data_print[31] vssd1 vssd1 vccd1 vccd1 _1137_/B sky130_fd_sc_hd__clkbuf_2
Xinput78 dout0_to_sram[3] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__buf_12
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput56 dout0_to_sram[12] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_8
Xinput67 dout0_to_sram[22] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_6
X_1556__663 vssd1 vssd1 vccd1 vccd1 _1556__663/HI la_data_out[4] sky130_fd_sc_hd__conb_1
Xinput89 la_data_in[13] vssd1 vssd1 vccd1 vccd1 _1693_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1516__A1 _2086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater657 _1767_/X vssd1 vssd1 vccd1 vccd1 _2149_/CLK sky130_fd_sc_hd__buf_12
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1225_ _1232_/A _1225_/B vssd1 vssd1 vccd1 vccd1 _1237_/B sky130_fd_sc_hd__or2_1
XFILLER_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1156_ _1148_/Y _1155_/X _1148_/Y _1155_/X vssd1 vssd1 vccd1 vccd1 _1156_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1087_ _2019_/Q _1087_/B vssd1 vssd1 vccd1 vccd1 _1088_/A sky130_fd_sc_hd__and2_1
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1989_ _1988_/X _1989_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1989_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1932__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input101_A la_data_in[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1443__B1 _2035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1994__A1 _1994_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2003__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1842__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0966__B _1721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output320_A _1887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1010_ _1010_/A vssd1 vssd1 vccd1 vccd1 _1010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2060__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1912_ _0906_/X _1912_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1912_/X sky130_fd_sc_hd__mux2_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1843_ _1842_/X input4/X _1942_/S vssd1 vssd1 vccd1 vccd1 _1843_/X sky130_fd_sc_hd__mux2_1
X_1774_ _1150_/A _1154_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1774_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1037__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1208_ _1208_/A _1221_/C vssd1 vssd1 vccd1 vccd1 _1208_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0892__A _1009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1139_ _2016_/X _1139_/B _2018_/Q vssd1 vssd1 vccd1 vccd1 _1140_/A sky130_fd_sc_hd__or3b_1
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1927__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput202 wr_data[118] vssd1 vssd1 vccd1 vccd1 _0972_/A sky130_fd_sc_hd__buf_2
Xinput235 wr_data[32] vssd1 vssd1 vccd1 vccd1 _1889_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input149_A la_data_in[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2083__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_49_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput213 wr_data[12] vssd1 vssd1 vccd1 vccd1 _1938_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput224 wr_data[22] vssd1 vssd1 vccd1 vccd1 _1978_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput257 wr_data[52] vssd1 vssd1 vccd1 vccd1 _1969_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput279 wr_data[72] vssd1 vssd1 vccd1 vccd1 _1920_/A1 sky130_fd_sc_hd__buf_2
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput268 wr_data[62] vssd1 vssd1 vccd1 vccd1 _2009_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput246 wr_data[42] vssd1 vssd1 vccd1 vccd1 _1929_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1416__B1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1837__S _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output368_A _1062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1490_ _2066_/Q _1486_/X input56/X _1487_/X vssd1 vssd1 vccd1 vccd1 _2066_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0977__A _0977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output535_A _2082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1668__775 vssd1 vssd1 vccd1 vccd1 _1668__775/HI la_data_out[117] sky130_fd_sc_hd__conb_1
XFILLER_121_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2111_ _1767_/X _2111_/D vssd1 vssd1 vccd1 vccd1 _2111_/Q sky130_fd_sc_hd__dfxtp_2
X_2042_ _2149_/CLK _2042_/D vssd1 vssd1 vccd1 vccd1 _2042_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1407__B1 input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1826_ _1825_/X _1689_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1826_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1757_ _1757_/A vssd1 vssd1 vccd1 vccd1 _1757_/X sky130_fd_sc_hd__buf_4
X_1688_ _1688_/A vssd1 vssd1 vccd1 vccd1 _1688_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0887__A _0887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1949__A1 _1949_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_126_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input266_A wr_data[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0990_ _0990_/A vssd1 vssd1 vccd1 vccd1 _0990_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output485_A _2037_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput517 _2066_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[44] sky130_fd_sc_hd__buf_2
Xoutput506 _2056_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[34] sky130_fd_sc_hd__buf_2
Xoutput539 _2086_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[64] sky130_fd_sc_hd__buf_2
XFILLER_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1542_ _2104_/Q _1540_/X input62/X _1541_/X vssd1 vssd1 vccd1 vccd1 _2104_/D sky130_fd_sc_hd__a22o_1
Xoutput528 _2076_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[54] sky130_fd_sc_hd__buf_2
XFILLER_113_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1473_ _1487_/A vssd1 vssd1 vccd1 vccd1 _1473_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1876__A0 _1336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2025_ _2155_/CLK _2025_/D vssd1 vssd1 vccd1 vccd1 _2025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1809_ _1209_/Y _1808_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1809_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1940__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__2121__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1398__A2 _1396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input77_A dout0_to_sram[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2011__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1135__B _1135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1858__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1850__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0974__B _1723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output400_A _1725_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_repeater648_A _1934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0973_ _0973_/A vssd1 vssd1 vccd1 vccd1 _0973_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_133_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput325 _1803_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[5] sky130_fd_sc_hd__buf_2
Xoutput314 _1851_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[13] sky130_fd_sc_hd__buf_2
XFILLER_99_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1525_ _2093_/Q _1519_/X input82/X _1520_/X vssd1 vssd1 vccd1 vccd1 _2093_/D sky130_fd_sc_hd__a22o_1
Xoutput369 _1064_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[26] sky130_fd_sc_hd__buf_2
Xoutput358 _1044_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[16] sky130_fd_sc_hd__buf_2
Xoutput347 _1687_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[7] sky130_fd_sc_hd__buf_2
Xoutput336 _1695_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[15] sky130_fd_sc_hd__buf_2
XFILLER_114_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1456_ input67/X _1452_/X _2044_/Q _1453_/X vssd1 vssd1 vccd1 vccd1 _2044_/D sky130_fd_sc_hd__o22a_1
XANTENNA__1045__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1387_ _2126_/Q _1382_/X input83/X _1383_/X vssd1 vssd1 vccd1 vccd1 _2126_/D sky130_fd_sc_hd__a22o_1
XANTENNA__2144__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1061__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2008_ _1006_/X _2008_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _2008_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1935__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input131_A la_data_in[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input229_A wr_data[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2006__S _2014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1845__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output350_A _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1146__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1310_ _1310_/A _1319_/B vssd1 vssd1 vccd1 vccd1 _1322_/B sky130_fd_sc_hd__or2_1
XANTENNA__0985__A _0985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output615_A _1076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1241_ _1244_/A _1239_/B _1240_/Y vssd1 vssd1 vccd1 vccd1 _1241_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1172_ input1/X _1150_/A _1168_/A _1168_/B vssd1 vssd1 vccd1 vccd1 _1173_/A sky130_fd_sc_hd__o211a_1
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0956_ _0956_/A _0972_/B vssd1 vssd1 vccd1 vccd1 _0957_/A sky130_fd_sc_hd__and2_1
XFILLER_137_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1231__A1 _1223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0887_ _0887_/A _1882_/S vssd1 vssd1 vccd1 vccd1 _0888_/A sky130_fd_sc_hd__and2_1
XANTENNA__0879__B _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1508_ _1508_/A vssd1 vssd1 vccd1 vccd1 _1508_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1439_ _1439_/A vssd1 vssd1 vccd1 vccd1 _1439_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0895__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1222__A1 _1210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input179_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_133_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output398_A _1723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1461__A1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 addr_in[2] vssd1 vssd1 vccd1 vccd1 _1168_/A sky130_fd_sc_hd__buf_2
X_1790_ _1789_/X _1683_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1790_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput46 core0_data_print[3] vssd1 vssd1 vccd1 vccd1 _1081_/B sky130_fd_sc_hd__buf_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput35 core0_data_print[22] vssd1 vssd1 vccd1 vccd1 _1119_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 core0_data_print[12] vssd1 vssd1 vccd1 vccd1 _1099_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_128_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput68 dout0_to_sram[23] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_8
XANTENNA_output565_A _2110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput79 dout0_to_sram[4] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__buf_8
Xinput57 dout0_to_sram[13] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_8
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1224_ _1228_/A vssd1 vssd1 vccd1 vccd1 _1232_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1155_ _0849_/Y _1151_/A _2152_/Q _1150_/A vssd1 vssd1 vccd1 vccd1 _1155_/X sky130_fd_sc_hd__o22a_1
XFILLER_37_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1086_ _1086_/A vssd1 vssd1 vccd1 vccd1 _1086_/X sky130_fd_sc_hd__buf_2
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1988_ _0986_/X _1988_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1988_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0939_ _0939_/A _0951_/B vssd1 vssd1 vccd1 vccd1 _0940_/A sky130_fd_sc_hd__and2_1
XFILLER_107_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_73_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1443__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input296_A wr_data[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1579__686 vssd1 vssd1 vccd1 vccd1 _1579__686/HI la_data_out[27] sky130_fd_sc_hd__conb_1
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_137_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_120_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_67_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_120_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1911_ _1910_/X _0900_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1911_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1434__A1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1842_ _1841_/X _1271_/Y _2013_/S vssd1 vssd1 vccd1 vccd1 _1842_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1773_ _1149_/Y _1772_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1773_/X sky130_fd_sc_hd__mux2_8
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1037__C _1747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1053__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1207_ _1204_/A _1196_/Y _1218_/B vssd1 vssd1 vccd1 vccd1 _1207_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1138_ _1138_/A vssd1 vssd1 vccd1 vccd1 _1138_/X sky130_fd_sc_hd__buf_2
XFILLER_41_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1069_ _1733_/A _2151_/Q _1763_/A vssd1 vssd1 vccd1 vccd1 _1070_/A sky130_fd_sc_hd__and3_1
XFILLER_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1943__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput203 wr_data[119] vssd1 vssd1 vccd1 vccd1 _0977_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1361__B1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput236 wr_data[33] vssd1 vssd1 vccd1 vccd1 _1893_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput225 wr_data[23] vssd1 vssd1 vccd1 vccd1 _1982_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput214 wr_data[13] vssd1 vssd1 vccd1 vccd1 _1942_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput258 wr_data[53] vssd1 vssd1 vccd1 vccd1 _1973_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput247 wr_data[43] vssd1 vssd1 vccd1 vccd1 _1933_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput269 wr_data[63] vssd1 vssd1 vccd1 vccd1 _2013_/A1 sky130_fd_sc_hd__buf_4
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input211_A wr_data[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input309_A wr_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1416__A1 _2147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2014__S _2014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1853__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0977__B _0993_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output528_A _2076_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output430_A _1983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2110_ _1767_/X _2110_/D vssd1 vssd1 vccd1 vccd1 _2110_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0993__A _0993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2041_ _2155_/CLK _2041_/D vssd1 vssd1 vccd1 vccd1 _2041_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1407__A1 _2140_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1825_ _1824_/X _1235_/A _1938_/S vssd1 vssd1 vccd1 vccd1 _1825_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1756_ _1756_/A vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1687_ _1687_/A vssd1 vssd1 vccd1 vccd1 _1687_/X sky130_fd_sc_hd__buf_4
XFILLER_131_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0887__B _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1894__A1 _1894_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1938__S _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2050__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_134_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input161_A la_data_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input259_A wr_data[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1885__A1 _1349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input22_A core0_data_print[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1702__A _1702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2009__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1848__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1594__701 vssd1 vssd1 vccd1 vccd1 _1594__701/HI la_data_out[42] sky130_fd_sc_hd__conb_1
XFILLER_13_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output380_A _1026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output478_A _2146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1635__742 vssd1 vssd1 vccd1 vccd1 _1635__742/HI la_data_out[83] sky130_fd_sc_hd__conb_1
Xoutput518 _2067_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[45] sky130_fd_sc_hd__buf_2
Xoutput507 _2057_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[35] sky130_fd_sc_hd__buf_2
X_1541_ _1541_/A vssd1 vssd1 vccd1 vccd1 _1541_/X sky130_fd_sc_hd__clkbuf_2
Xoutput529 _2077_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[55] sky130_fd_sc_hd__buf_2
XANTENNA_output645_A _1092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1472_ _1508_/A vssd1 vssd1 vccd1 vccd1 _1487_/A sky130_fd_sc_hd__buf_2
XFILLER_113_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_2024_ _2155_/CLK _2024_/D vssd1 vssd1 vccd1 vccd1 _2024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2073__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1059__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1808_ _1807_/X _1686_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1808_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0898__A _0898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1739_ _1739_/A vssd1 vssd1 vccd1 vccd1 _1739_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1867__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1619__726 vssd1 vssd1 vccd1 vccd1 _1619__726/HI la_data_out[67] sky130_fd_sc_hd__conb_1
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1432__A _1439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2096__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output595_A _1757_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0972_ _0972_/A _0972_/B vssd1 vssd1 vccd1 vccd1 _0973_/A sky130_fd_sc_hd__and2_1
XFILLER_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput315 _1857_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[14] sky130_fd_sc_hd__buf_2
Xoutput326 _1809_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[6] sky130_fd_sc_hd__buf_2
Xoutput337 _1696_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[16] sky130_fd_sc_hd__buf_2
Xoutput348 _1688_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[8] sky130_fd_sc_hd__buf_2
XANTENNA__1546__B1 input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1524_ _2092_/Q _1519_/X input81/X _1520_/X vssd1 vssd1 vccd1 vccd1 _2092_/D sky130_fd_sc_hd__a22o_1
Xoutput359 _1046_/X vssd1 vssd1 vccd1 vccd1 data_out_to_core[17] sky130_fd_sc_hd__buf_2
XFILLER_5_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1455_ input66/X _1452_/X _2043_/Q _1453_/X vssd1 vssd1 vccd1 vccd1 _2043_/D sky130_fd_sc_hd__o22a_1
XFILLER_68_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1386_ _2125_/Q _1382_/X input82/X _1383_/X vssd1 vssd1 vccd1 vccd1 _2125_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1045__C _1751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1849__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2007_ _2006_/X _1000_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _2007_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1061__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1537__B1 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1951__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input124_A la_data_in[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1528__B1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output343_A _1683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1861__S _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0985__B _0993_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1240_ _1250_/B vssd1 vssd1 vccd1 vccd1 _1240_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output510_A _2060_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1171_ _1175_/B _1170_/B _1182_/B vssd1 vssd1 vccd1 vccd1 _1171_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA_output608_A _1740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2008__A1 _2008_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0955_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0972_/B sky130_fd_sc_hd__clkbuf_4
X_0886_ _0886_/A vssd1 vssd1 vccd1 vccd1 _0886_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2111__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1507_ _1507_/A vssd1 vssd1 vccd1 vccd1 _1507_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1771__S _1922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1438_ _1438_/A vssd1 vssd1 vccd1 vccd1 _1438_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0895__B _1704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1369_ _2117_/Q _1366_/X input77/X _1367_/X vssd1 vssd1 vccd1 vccd1 _2117_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1946__S _2010_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_127_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1930__A0 _1929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input241_A wr_data[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1710__A _1710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2134__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1856__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput25 core0_data_print[13] vssd1 vssd1 vccd1 vccd1 _1101_/B sky130_fd_sc_hd__buf_2
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput36 core0_data_print[23] vssd1 vssd1 vccd1 vccd1 _1121_/B sky130_fd_sc_hd__clkbuf_2
Xinput14 addr_in[3] vssd1 vssd1 vccd1 vccd1 _1168_/B sky130_fd_sc_hd__clkbuf_2
Xinput58 dout0_to_sram[14] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_8
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput47 core0_data_print[4] vssd1 vssd1 vccd1 vccd1 _1083_/B sky130_fd_sc_hd__buf_2
XANTENNA_output460_A _2130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput69 dout0_to_sram[24] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_6
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_109_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1921__A0 _1920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1223_ _1223_/A vssd1 vssd1 vccd1 vccd1 _1228_/A sky130_fd_sc_hd__inv_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater648 _1934_/S vssd1 vssd1 vccd1 vccd1 _2014_/S sky130_fd_sc_hd__buf_4
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1154_ _1154_/A vssd1 vssd1 vccd1 vccd1 _1154_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1085_ _2019_/Q _1085_/B vssd1 vssd1 vccd1 vccd1 _1086_/A sky130_fd_sc_hd__and2_1
XFILLER_21_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1987_ _1986_/X _0980_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1987_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0938_ _0938_/A vssd1 vssd1 vccd1 vccd1 _0938_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1067__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0869_ _2155_/Q vssd1 vssd1 vccd1 vccd1 _0870_/A sky130_fd_sc_hd__inv_2
XFILLER_130_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_113_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input191_A wr_data[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input289_A wr_data[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input52_A core0_data_print[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1705__A _1705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ _1909_/X _1910_/A1 _1938_/S vssd1 vssd1 vccd1 vccd1 _1910_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ _1840_/X _1273_/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1841_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1772_ _1771_/X _1680_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1772_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__C _1755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1206_ _1208_/A _1206_/B vssd1 vssd1 vccd1 vccd1 _1218_/B sky130_fd_sc_hd__or2_1
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1137_ _2019_/Q _1137_/B vssd1 vssd1 vccd1 vccd1 _1138_/A sky130_fd_sc_hd__and2_1
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1068_ _1068_/A vssd1 vssd1 vccd1 vccd1 _1068_/X sky130_fd_sc_hd__buf_4
XFILLER_41_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1652__759 vssd1 vssd1 vccd1 vccd1 _1652__759/HI la_data_out[101] sky130_fd_sc_hd__conb_1
XFILLER_134_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1361__A1 _2111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput226 wr_data[24] vssd1 vssd1 vccd1 vccd1 _1986_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput204 wr_data[11] vssd1 vssd1 vccd1 vccd1 _1934_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput215 wr_data[14] vssd1 vssd1 vccd1 vccd1 _1946_/A1 sky130_fd_sc_hd__buf_4
Xinput237 wr_data[34] vssd1 vssd1 vccd1 vccd1 _1897_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput259 wr_data[54] vssd1 vssd1 vccd1 vccd1 _1977_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput248 wr_data[44] vssd1 vssd1 vccd1 vccd1 _1937_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input204_A wr_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1352__A1 _1349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2040_ _2155_/CLK _2040_/D vssd1 vssd1 vccd1 vccd1 _2040_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0993__B _0993_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1824_ _1823_/X _1238_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1824_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1755_ _1755_/A vssd1 vssd1 vccd1 vccd1 _1755_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1686_ _1686_/A vssd1 vssd1 vccd1 vccd1 _1686_/X sky130_fd_sc_hd__buf_2
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1954__S _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input154_A la_data_in[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input15_A addr_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_138_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1674__781 vssd1 vssd1 vccd1 vccd1 _1674__781/HI la_data_out[123] sky130_fd_sc_hd__conb_1
X_1540_ _1540_/A vssd1 vssd1 vccd1 vccd1 _1540_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput508 _2058_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[36] sky130_fd_sc_hd__buf_2
XANTENNA__1864__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput519 _2068_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[46] sky130_fd_sc_hd__buf_2
XFILLER_114_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_114_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output638_A _1136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1471_ _1507_/A vssd1 vssd1 vccd1 vccd1 _1508_/A sky130_fd_sc_hd__inv_2
XANTENNA_output540_A _2087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2023_ _2155_/CLK _2023_/D vssd1 vssd1 vccd1 vccd1 _2023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1059__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1807_ _1806_/X _1204_/A _1922_/S vssd1 vssd1 vccd1 vccd1 _1807_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1774__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1738_ _1738_/A vssd1 vssd1 vccd1 vccd1 _1738_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1075__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A addr_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1949__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1658__765 vssd1 vssd1 vccd1 vccd1 _1658__765/HI la_data_out[107] sky130_fd_sc_hd__conb_1
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input271_A wr_data[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1713__A _1713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1859__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1491__B1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ _0971_/A vssd1 vssd1 vccd1 vccd1 _0971_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output588_A _1751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0999__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput316 _1863_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[15] sky130_fd_sc_hd__buf_2
Xoutput327 _1815_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[7] sky130_fd_sc_hd__buf_2
XFILLER_126_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1523_ _2091_/Q _1519_/X input80/X _1520_/X vssd1 vssd1 vccd1 vccd1 _2091_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput338 _1697_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[17] sky130_fd_sc_hd__buf_2
Xoutput349 _1689_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[9] sky130_fd_sc_hd__buf_2
XFILLER_114_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1454_ input65/X _1452_/X _2042_/Q _1453_/X vssd1 vssd1 vccd1 vccd1 _2042_/D sky130_fd_sc_hd__o22a_1
XFILLER_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1385_ _2124_/Q _1382_/X input81/X _1383_/X vssd1 vssd1 vccd1 vccd1 _2124_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2006_ _2005_/X _2006_/A1 _2014_/S vssd1 vssd1 vccd1 vccd1 _2006_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1061__C _1759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2040__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1769__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1482__B1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1537__A1 _2101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1537__B2 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input117_A la_data_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input82_A dout0_to_sram[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1708__A _1708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1528__A1 _2094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_110_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2063__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1170_ _1175_/B _1170_/B vssd1 vssd1 vccd1 vccd1 _1182_/B sky130_fd_sc_hd__or2_1
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output503_A _2053_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1464__B1 _2050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater653_A _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0954_ _0954_/A vssd1 vssd1 vccd1 vccd1 _0954_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1767__A1 _1767_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0885_ _1732_/A _1702_/A vssd1 vssd1 vccd1 vccd1 _0886_/A sky130_fd_sc_hd__and2_1
XFILLER_119_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1506_ _2078_/Q _1500_/X input69/X _1501_/X vssd1 vssd1 vccd1 vccd1 _2078_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1437_ input84/X _1431_/X _2031_/Q _1432_/X vssd1 vssd1 vccd1 vccd1 _2031_/D sky130_fd_sc_hd__o22a_1
X_1368_ _2116_/Q _1366_/X input76/X _1367_/X vssd1 vssd1 vccd1 vccd1 _2116_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1299_ _1302_/A _1310_/A vssd1 vssd1 vccd1 vccd1 _1299_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1455__B1 _2043_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1962__S _1990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2086__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input234_A wr_data[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput37 core0_data_print[24] vssd1 vssd1 vccd1 vccd1 _1123_/B sky130_fd_sc_hd__clkbuf_4
Xinput15 addr_in[4] vssd1 vssd1 vccd1 vccd1 _1177_/A sky130_fd_sc_hd__buf_6
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 core0_data_print[14] vssd1 vssd1 vccd1 vccd1 _1103_/B sky130_fd_sc_hd__buf_2
XANTENNA__1438__A _1438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput59 dout0_to_sram[15] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_6
Xinput48 core0_data_print[5] vssd1 vssd1 vccd1 vccd1 _1085_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output453_A _2123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1872__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output620_A _1104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1222_ _1210_/A _1208_/Y _1232_/B vssd1 vssd1 vccd1 vccd1 _1222_/X sky130_fd_sc_hd__o21a_1
Xrepeater649 _1942_/S vssd1 vssd1 vccd1 vccd1 _1934_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1153_ _1144_/X _1160_/A _1168_/C vssd1 vssd1 vccd1 vccd1 _1154_/A sky130_fd_sc_hd__a21oi_1
XFILLER_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1084_ _1084_/A vssd1 vssd1 vccd1 vccd1 _1084_/X sky130_fd_sc_hd__buf_2
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1988__A1 _1988_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1986_ _1985_/X _1986_/A1 _1990_/S vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0937_ _1732_/A _1714_/A vssd1 vssd1 vccd1 vccd1 _0938_/A sky130_fd_sc_hd__and2_1
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1067__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0868_ _0868_/A vssd1 vssd1 vccd1 vccd1 _2015_/S sky130_fd_sc_hd__buf_12
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1782__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1912__A1 _1912_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1083__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1957__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input184_A wr_data[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input45_A core0_data_print[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1721__A _1721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2101__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1867__S _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1840_ input4/X _1276_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1840_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output570_A _2114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1771_ _1770_/X input1/X _1922_/S vssd1 vssd1 vccd1 vccd1 _1771_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1205_ _1204_/A _1204_/B _1215_/B vssd1 vssd1 vccd1 vccd1 _1205_/X sky130_fd_sc_hd__o21a_1
X_1136_ _1136_/A vssd1 vssd1 vccd1 vccd1 _1136_/X sky130_fd_sc_hd__buf_2
XFILLER_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_25_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1067_ _1733_/A _2151_/Q _1762_/A vssd1 vssd1 vccd1 vccd1 _1068_/A sky130_fd_sc_hd__and3_1
XFILLER_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1777__S _1922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1969_ _1968_/X _1969_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1969_/X sky130_fd_sc_hd__mux2_2
XFILLER_135_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput205 wr_data[120] vssd1 vssd1 vccd1 vccd1 _0981_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput227 wr_data[25] vssd1 vssd1 vccd1 vccd1 _1990_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput216 wr_data[15] vssd1 vssd1 vccd1 vccd1 _1950_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput249 wr_data[45] vssd1 vssd1 vccd1 vccd1 _1941_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput238 wr_data[35] vssd1 vssd1 vccd1 vccd1 _1901_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2124__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1585__692 vssd1 vssd1 vccd1 vccd1 _1585__692/HI la_data_out[33] sky130_fd_sc_hd__conb_1
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_125_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1716__A _1716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_117_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1823_ _1822_/X _1241_/Y _2012_/S vssd1 vssd1 vccd1 vccd1 _1823_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1754_ _1754_/A vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1685_ _1685_/A vssd1 vssd1 vccd1 vccd1 _1685_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2147__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1569__676 vssd1 vssd1 vccd1 vccd1 _1569__676/HI la_data_out[17] sky130_fd_sc_hd__conb_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2099_ _1767_/X _2099_/D vssd1 vssd1 vccd1 vccd1 _2099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1119_ _2019_/Q _1119_/B vssd1 vssd1 vccd1 vccd1 _1120_/A sky130_fd_sc_hd__and2_1
XFILLER_110_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_123_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1970__S _2014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input147_A la_data_in[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput509 _2059_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[37] sky130_fd_sc_hd__buf_2
XFILLER_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1470_ _1486_/A vssd1 vssd1 vccd1 vccd1 _1470_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output533_A _2081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1880__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2022_ _2155_/CLK _2022_/D vssd1 vssd1 vccd1 vccd1 _2022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1059__C _1758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1806_ _1805_/X _1203_/Y _2013_/S vssd1 vssd1 vccd1 vccd1 _1806_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1737_ _1737_/A vssd1 vssd1 vccd1 vccd1 _1737_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1075__B _1075_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1790__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1091__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1965__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input264_A wr_data[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0970_ _1732_/A _1722_/A vssd1 vssd1 vccd1 vccd1 _0971_/A sky130_fd_sc_hd__and2_1
XFILLER_60_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output483_A _2035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1875__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0999__B _1729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput317 _1869_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[16] sky130_fd_sc_hd__buf_2
Xoutput339 _1698_/X vssd1 vssd1 vccd1 vccd1 addr_to_core_mem[18] sky130_fd_sc_hd__buf_2
XFILLER_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1522_ _2090_/Q _1519_/X input79/X _1520_/X vssd1 vssd1 vccd1 vccd1 _2090_/D sky130_fd_sc_hd__a22o_1
Xoutput328 _1821_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[8] sky130_fd_sc_hd__buf_2
XFILLER_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1453_ _1460_/A vssd1 vssd1 vccd1 vccd1 _1453_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1384_ _2123_/Q _1382_/X input80/X _1383_/X vssd1 vssd1 vccd1 vccd1 _2123_/D sky130_fd_sc_hd__a22o_1
XFILLER_95_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2005_ _2004_/X _2005_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _2005_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_36_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1482__A1 _2060_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1785__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1537__A2 _1533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_120_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1625__732 vssd1 vssd1 vccd1 vccd1 _1625__732/HI la_data_out[73] sky130_fd_sc_hd__conb_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input75_A dout0_to_sram[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1724__A _1724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output329_A _1827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1464__A1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0953_ _1732_/A _1718_/A vssd1 vssd1 vccd1 vccd1 _0954_/A sky130_fd_sc_hd__and2_1
X_0884_ _0884_/A vssd1 vssd1 vccd1 vccd1 _0884_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1505_ _2077_/Q _1500_/X input68/X _1501_/X vssd1 vssd1 vccd1 vccd1 _2077_/D sky130_fd_sc_hd__a22o_1
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1436_ input83/X _1431_/X _2030_/Q _1432_/X vssd1 vssd1 vccd1 vccd1 _2030_/D sky130_fd_sc_hd__o22a_1
XFILLER_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1367_ _1520_/A vssd1 vssd1 vccd1 vccd1 _1367_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1609__716 vssd1 vssd1 vccd1 vccd1 _1609__716/HI la_data_out[57] sky130_fd_sc_hd__conb_1
XFILLER_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1298_ _1297_/A _1308_/A _1297_/Y vssd1 vssd1 vccd1 vccd1 _1298_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1455__B2 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1455__A1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1391__B1 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input227_A wr_data[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1719__A _1719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 addr_in[5] vssd1 vssd1 vccd1 vccd1 _1189_/A sky130_fd_sc_hd__buf_4
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput27 core0_data_print[15] vssd1 vssd1 vccd1 vccd1 _1105_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_109_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput49 core0_data_print[6] vssd1 vssd1 vccd1 vccd1 _1087_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 core0_data_print[25] vssd1 vssd1 vccd1 vccd1 _1125_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2030__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output446_A _1927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1221_ _1221_/A _1221_/B _1221_/C vssd1 vssd1 vccd1 vccd1 _1232_/B sky130_fd_sc_hd__or3_1
XFILLER_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1152_ _1152_/A _1160_/A vssd1 vssd1 vccd1 vccd1 _1168_/C sky130_fd_sc_hd__nor2_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1083_ _2019_/Q _1083_/B vssd1 vssd1 vccd1 vccd1 _1084_/A sky130_fd_sc_hd__and2_1
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1437__A1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ _1984_/X _1985_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1985_/X sky130_fd_sc_hd__mux2_1
X_0936_ _0936_/A vssd1 vssd1 vccd1 vccd1 _0936_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1067__C _1762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0867_ _0867_/A _1732_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _0868_/A sky130_fd_sc_hd__or3b_1
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1083__B _1083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1419_ _1419_/A vssd1 vssd1 vccd1 vccd1 _2019_/D sky130_fd_sc_hd__clkinv_2
XFILLER_130_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1428__A1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1428__B2 _1425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2053__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1973__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input177_A requested vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1364__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input38_A core0_data_print[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output396_A _1721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1770_ _1769_/X _1144_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1770_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1883__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1204_ _1204_/A _1204_/B vssd1 vssd1 vccd1 vccd1 _1215_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1135_ _2019_/Q _1135_/B vssd1 vssd1 vccd1 vccd1 _1136_/A sky130_fd_sc_hd__and2_1
XFILLER_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1066_ _1066_/A vssd1 vssd1 vccd1 vccd1 _1066_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2076__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_119_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1968_ _0965_/X _1968_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1968_/X sky130_fd_sc_hd__mux2_2
X_1899_ _1898_/X _0886_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1899_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0919_ _0919_/A vssd1 vssd1 vccd1 vccd1 _0919_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1793__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput206 wr_data[121] vssd1 vssd1 vccd1 vccd1 _0985_/A sky130_fd_sc_hd__buf_2
XFILLER_130_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput217 wr_data[16] vssd1 vssd1 vccd1 vccd1 _1954_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput239 wr_data[36] vssd1 vssd1 vccd1 vccd1 _1905_/A1 sky130_fd_sc_hd__buf_2
Xinput228 wr_data[26] vssd1 vssd1 vccd1 vccd1 _1994_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1968__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input294_A wr_data[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_125_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0901__A _0901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1732__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output311_A _1833_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2099__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1878__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1822_ _1235_/A _1243_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1822_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1753_ _1753_/A vssd1 vssd1 vccd1 vccd1 _1753_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1684_ _1684_/A vssd1 vssd1 vccd1 vccd1 _1684_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1879__A1 _1336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ _2149_/CLK _2098_/D vssd1 vssd1 vccd1 vccd1 _2098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1118_ _1118_/A vssd1 vssd1 vccd1 vccd1 _1118_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1788__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1049_ _1733_/A _2151_/Q _1753_/A vssd1 vssd1 vccd1 vccd1 _1050_/A sky130_fd_sc_hd__and3_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1089__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_130_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input307_A wr_data[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1727__A _1727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_95_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output526_A _2074_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2021_ _2155_/CLK _2152_/Q vssd1 vssd1 vccd1 vccd1 _2021_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1642__749 vssd1 vssd1 vccd1 vccd1 _1642__749/HI la_data_out[90] sky130_fd_sc_hd__conb_1
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2114__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1805_ _1804_/X _1205_/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1805_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1736_ _1736_/A vssd1 vssd1 vccd1 vccd1 _1736_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1091__B _1091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1981__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input257_A wr_data[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input20_A addr_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2137__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output476_A _2144_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1521_ _2089_/Q _1519_/X input78/X _1520_/X vssd1 vssd1 vccd1 vccd1 _2089_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1891__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput318 _1875_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[17] sky130_fd_sc_hd__buf_2
XFILLER_5_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput329 _1827_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[9] sky130_fd_sc_hd__buf_2
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1452_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1452_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1383_ _1390_/A vssd1 vssd1 vccd1 vccd1 _1383_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2004_ _1002_/X _2004_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _2004_/X sky130_fd_sc_hd__mux2_2
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1719_ _1719_/A vssd1 vssd1 vccd1 vccd1 _1719_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1942__A0 _1941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1664__771 vssd1 vssd1 vccd1 vccd1 _1664__771/HI la_data_out[113] sky130_fd_sc_hd__conb_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1976__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input68_A dout0_to_sram[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1161__A1 _1150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1740__A _1740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1886__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0952_ _0952_/A vssd1 vssd1 vccd1 vccd1 _0952_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0883_ _0883_/A _1882_/S vssd1 vssd1 vccd1 vccd1 _0884_/A sky130_fd_sc_hd__and2_1
XFILLER_133_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1504_ _2076_/Q _1500_/X input67/X _1501_/X vssd1 vssd1 vccd1 vccd1 _2076_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1924__A0 _0919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1435_ input82/X _1431_/X _2029_/Q _1432_/X vssd1 vssd1 vccd1 vccd1 _2029_/D sky130_fd_sc_hd__o22a_1
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1366_ _1519_/A vssd1 vssd1 vccd1 vccd1 _1366_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1648__755 vssd1 vssd1 vccd1 vccd1 _1648__755/HI la_data_out[96] sky130_fd_sc_hd__conb_1
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1297_ _1297_/A _1308_/A vssd1 vssd1 vccd1 vccd1 _1297_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1455__A2 _1452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1796__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1097__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input122_A la_data_in[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput28 core0_data_print[16] vssd1 vssd1 vccd1 vccd1 _1107_/B sky130_fd_sc_hd__buf_2
Xinput17 addr_in[6] vssd1 vssd1 vccd1 vccd1 _1204_/A sky130_fd_sc_hd__buf_2
Xinput39 core0_data_print[26] vssd1 vssd1 vccd1 vccd1 _1127_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1735__A _1735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1906__A0 _1905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1220_ _1218_/A _1218_/B _1219_/Y vssd1 vssd1 vccd1 vccd1 _1220_/Y sky130_fd_sc_hd__a21oi_1
X_1151_ _1151_/A vssd1 vssd1 vccd1 vccd1 _1160_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output606_A _1738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1082_ _1082_/A vssd1 vssd1 vccd1 vccd1 _1082_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1984_ _0982_/X _1984_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1984_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0935_ _0935_/A _0951_/B vssd1 vssd1 vccd1 vccd1 _0936_/A sky130_fd_sc_hd__and2_1
XFILLER_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0866_ _0866_/A vssd1 vssd1 vccd1 vccd1 _0867_/A sky130_fd_sc_hd__inv_2
XFILLER_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1418_ _2149_/Q _1389_/A input77/X _1390_/A vssd1 vssd1 vccd1 vccd1 _2149_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1349_ _1349_/A vssd1 vssd1 vccd1 vccd1 _1349_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1428__A2 _1422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_4_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1364__A1 _2114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput490 _2023_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output389_A _1715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output556_A _2029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1203_ _1208_/A _1202_/B _1202_/Y vssd1 vssd1 vccd1 vccd1 _1203_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1134_ _1134_/A vssd1 vssd1 vccd1 vccd1 _1134_/X sky130_fd_sc_hd__buf_2
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1065_ _1733_/A _2151_/Q _1761_/A vssd1 vssd1 vccd1 vccd1 _1066_/A sky130_fd_sc_hd__and3_1
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1967_ _1966_/X _0959_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1967_/X sky130_fd_sc_hd__mux2_2
X_1898_ _1897_/X _1898_/A1 _1934_/S vssd1 vssd1 vccd1 vccd1 _1898_/X sky130_fd_sc_hd__mux2_1
X_0918_ _0918_/A _0930_/B vssd1 vssd1 vccd1 vccd1 _0919_/A sky130_fd_sc_hd__and2_2
XFILLER_107_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0849_ _2152_/Q vssd1 vssd1 vccd1 vccd1 _0849_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput207 wr_data[122] vssd1 vssd1 vccd1 vccd1 _0989_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput218 wr_data[17] vssd1 vssd1 vccd1 vccd1 _1958_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput229 wr_data[27] vssd1 vssd1 vccd1 vccd1 _1998_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2020__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1984__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input287_A wr_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0901__B _0909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input50_A core0_data_print[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1821_ _1234_/Y _1820_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1821_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1894__S _1990_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1752_ _1752_/A vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1683_ _1683_/A vssd1 vssd1 vccd1 vccd1 _1683_/X sky130_fd_sc_hd__buf_4
XANTENNA__1328__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2043__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1117_ _2019_/Q _1117_/B vssd1 vssd1 vccd1 vccd1 _1118_/A sky130_fd_sc_hd__and2_1
X_2097_ _2149_/CLK _2097_/D vssd1 vssd1 vccd1 vccd1 _2097_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1048_ _1048_/A vssd1 vssd1 vccd1 vccd1 _1048_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1089__B _1089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1979__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input202_A wr_data[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input98_A la_data_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2066__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output421_A _1951_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output519_A _2068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2020_ _2155_/CLK _2154_/Q vssd1 vssd1 vccd1 vccd1 _2020_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__1889__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_51_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1804_ _1204_/A _1207_/X _1882_/S vssd1 vssd1 vccd1 vccd1 _1804_/X sky130_fd_sc_hd__mux2_1
X_1735_ _1735_/A vssd1 vssd1 vccd1 vccd1 _1735_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1575__682 vssd1 vssd1 vccd1 vccd1 _1575__682/HI la_data_out[23] sky130_fd_sc_hd__conb_1
XFILLER_104_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1799__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2149_ _2149_/CLK _2149_/D vssd1 vssd1 vccd1 vccd1 _2149_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__1485__B1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_135_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_5_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2089__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input152_A la_data_in[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0907__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1476__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A addr_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1738__A _1738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1559__666 vssd1 vssd1 vccd1 vccd1 _1559__666/HI la_data_out[7] sky130_fd_sc_hd__conb_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output371_A _1068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output469_A _2138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1520_ _1520_/A vssd1 vssd1 vccd1 vccd1 _1520_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput319 _1881_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[18] sky130_fd_sc_hd__buf_2
XANTENNA__1400__B1 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output636_A _1134_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1451_ input63/X _1445_/X _2041_/Q _1446_/X vssd1 vssd1 vccd1 vccd1 _2041_/D sky130_fd_sc_hd__o22a_1
XFILLER_4_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1382_ _1389_/A vssd1 vssd1 vccd1 vccd1 _1382_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1473__A _1487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1467__B1 _2053_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2003_ _2002_/X _0996_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _2003_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1718_ _1718_/A vssd1 vssd1 vccd1 vccd1 _1718_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1942__A1 _1942_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A addr_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1458__B1 _2046_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1992__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2104__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1449__B1 _2039_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0951_ _0951_/A _0951_/B vssd1 vssd1 vccd1 vccd1 _0952_/A sky130_fd_sc_hd__and2_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1468__A _2021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output586_A _1749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0882_ _0882_/A vssd1 vssd1 vccd1 vccd1 _0882_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1503_ _2075_/Q _1500_/X input66/X _1501_/X vssd1 vssd1 vccd1 vccd1 _2075_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1434_ input81/X _1431_/X _2028_/Q _1432_/X vssd1 vssd1 vccd1 vccd1 _2028_/D sky130_fd_sc_hd__o22a_1
X_1365_ _2115_/Q _1357_/X input74/X _1360_/X vssd1 vssd1 vccd1 vccd1 _2115_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1296_ input6/X _1285_/Y _1305_/B vssd1 vssd1 vccd1 vccd1 _1296_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2127__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input115_A la_data_in[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1987__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input80_A dout0_to_sram[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 addr_in[7] vssd1 vssd1 vccd1 vccd1 _1210_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_109_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput29 core0_data_print[17] vssd1 vssd1 vccd1 vccd1 _1109_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_136_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0920__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1751__A _1751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1150_ _1150_/A vssd1 vssd1 vccd1 vccd1 _1151_/A sky130_fd_sc_hd__inv_2
XFILLER_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1081_ _2019_/Q _1081_/B vssd1 vssd1 vccd1 vccd1 _1082_/A sky130_fd_sc_hd__and2_1
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1897__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_repeater651_A _1954_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ _1982_/X _0975_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1983_/X sky130_fd_sc_hd__mux2_2
X_0934_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0951_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0865_ _0865_/A vssd1 vssd1 vccd1 vccd1 _0865_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1615__722 vssd1 vssd1 vccd1 vccd1 _1615__722/HI la_data_out[63] sky130_fd_sc_hd__conb_1
XFILLER_88_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1417_ _2148_/Q _1389_/A input76/X _1390_/A vssd1 vssd1 vccd1 vccd1 _2148_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_84_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1348_ _1341_/A _1346_/B _1347_/Y vssd1 vssd1 vccd1 vccd1 _1348_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1279_ _1274_/A _1277_/B _1278_/Y vssd1 vssd1 vccd1 vccd1 _1279_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2010__A0 _2009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput480 _2148_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[126] sky130_fd_sc_hd__buf_2
Xoutput491 _2042_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input232_A wr_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1746__A _1746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output549_A _2095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1202_ _1208_/A _1202_/B vssd1 vssd1 vccd1 vccd1 _1202_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_93_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1133_ _2019_/Q _1133_/B vssd1 vssd1 vccd1 vccd1 _1134_/A sky130_fd_sc_hd__and2_1
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1064_ _1064_/A vssd1 vssd1 vccd1 vccd1 _1064_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1966_ _1965_/X _1966_/A1 _2010_/S vssd1 vssd1 vccd1 vccd1 _1966_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0917_ _0917_/A vssd1 vssd1 vccd1 vccd1 _0917_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1897_ _1896_/X _1897_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1897_/X sky130_fd_sc_hd__mux2_2
XFILLER_134_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0848_ _1148_/A vssd1 vssd1 vccd1 vccd1 _0875_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput208 wr_data[123] vssd1 vssd1 vccd1 vccd1 _0993_/A sky130_fd_sc_hd__buf_4
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_130_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput219 wr_data[18] vssd1 vssd1 vccd1 vccd1 _1962_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input182_A wr_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1592__699 vssd1 vssd1 vccd1 vccd1 _1592__699/HI la_data_out[40] sky130_fd_sc_hd__conb_1
XFILLER_106_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input43_A core0_data_print[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1273__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output499_A _2050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1820_ _1819_/X _1688_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1820_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1751_ _1751_/A vssd1 vssd1 vccd1 vccd1 _1751_/X sky130_fd_sc_hd__buf_4
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1682_ _1682_/A vssd1 vssd1 vccd1 vccd1 _1682_/X sky130_fd_sc_hd__buf_4
XFILLER_132_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1116_ _1116_/A vssd1 vssd1 vccd1 vccd1 _1116_/X sky130_fd_sc_hd__clkbuf_2
X_2096_ _2149_/CLK _2096_/D vssd1 vssd1 vccd1 vccd1 _2096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1047_ _1733_/A _2151_/Q _1752_/A vssd1 vssd1 vccd1 vccd1 _1048_/A sky130_fd_sc_hd__and3_1
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1264__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1949_ _1948_/X _1949_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1949_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1995__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output414_A _1709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1803_ _1199_/X _1802_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1803_/X sky130_fd_sc_hd__mux2_4
XFILLER_129_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1734_ _1734_/A vssd1 vssd1 vccd1 vccd1 _1734_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2148_ _1767_/X _2148_/D vssd1 vssd1 vccd1 vccd1 _2148_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__1485__A1 _2063_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2079_ _1767_/X _2079_/D vssd1 vssd1 vccd1 vccd1 _2079_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_108_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input145_A la_data_in[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1476__B2 _1473_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1476__A1 _2056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2033__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1400__A1 _2135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1754__A _1754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output364_A _1054_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1400__B2 _1397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1450_ input62/X _1445_/X _2040_/Q _1446_/X vssd1 vssd1 vccd1 vccd1 _2040_/D sky130_fd_sc_hd__o22a_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1381_ _2122_/Q _1373_/X input79/X _1376_/X vssd1 vssd1 vccd1 vccd1 _2122_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output531_A _2079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output629_A _1120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1467__A1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1467__B2 _1439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2002_ _2001_/X _2002_/A1 _2010_/S vssd1 vssd1 vccd1 vccd1 _2002_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1717_ _1717_/A vssd1 vssd1 vccd1 vccd1 _1717_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1155__B1 _2152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1458__B2 _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1458__A1 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2056__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1394__B1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1632__739 vssd1 vssd1 vccd1 vccd1 _1632__739/HI la_data_out[80] sky130_fd_sc_hd__conb_1
XFILLER_123_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input262_A wr_data[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1449__A1 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0950_ _0950_/A vssd1 vssd1 vccd1 vccd1 _0950_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1749__A _1749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output481_A _2149_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0881_ _1732_/A _1701_/A vssd1 vssd1 vccd1 vccd1 _0882_/A sky130_fd_sc_hd__and2_1
XFILLER_9_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1385__B1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_126_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1502_ _2074_/Q _1500_/X input65/X _1501_/X vssd1 vssd1 vccd1 vccd1 _2074_/D sky130_fd_sc_hd__a22o_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1433_ input80/X _1431_/X _2027_/Q _1432_/X vssd1 vssd1 vccd1 vccd1 _2027_/D sky130_fd_sc_hd__o22a_1
X_1364_ _2114_/Q _1357_/X input73/X _1360_/X vssd1 vssd1 vccd1 vccd1 _2114_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_110_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1295_ _1302_/A _1295_/B vssd1 vssd1 vccd1 vccd1 _1305_/B sky130_fd_sc_hd__or2_1
XFILLER_49_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2079__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput640 _1082_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input108_A la_data_in[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput19 addr_in[8] vssd1 vssd1 vccd1 vccd1 _1223_/A sky130_fd_sc_hd__buf_4
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input73_A dout0_to_sram[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0920__B _1710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output327_A _1815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1080_ _1080_/A vssd1 vssd1 vccd1 vccd1 _1080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ _1981_/X _1982_/A1 _2010_/S vssd1 vssd1 vccd1 vccd1 _1982_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0933_ _0933_/A vssd1 vssd1 vccd1 vccd1 _0933_/X sky130_fd_sc_hd__clkbuf_1
X_0864_ _1700_/A _1732_/A vssd1 vssd1 vccd1 vccd1 _0865_/A sky130_fd_sc_hd__and2_1
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1654__761 vssd1 vssd1 vccd1 vccd1 _1654__761/HI la_data_out[103] sky130_fd_sc_hd__conb_1
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1416_ _2147_/Q _1410_/X input74/X _1411_/X vssd1 vssd1 vccd1 vccd1 _2147_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1347_ _1347_/A vssd1 vssd1 vccd1 vccd1 _1347_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1530__B1 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1278_ _1289_/B vssd1 vssd1 vccd1 vccd1 _1278_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2010__A1 _2010_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput470 _2139_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[117] sky130_fd_sc_hd__buf_2
XFILLER_106_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput481 _2149_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[127] sky130_fd_sc_hd__buf_2
Xoutput492 _2043_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[21] sky130_fd_sc_hd__buf_2
XFILLER_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1521__B1 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1998__S _2014_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input225_A wr_data[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1597__704 vssd1 vssd1 vccd1 vccd1 _1597__704/HI la_data_out[45] sky130_fd_sc_hd__conb_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0931__A _0931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1638__745 vssd1 vssd1 vccd1 vccd1 _1638__745/HI la_data_out[86] sky130_fd_sc_hd__conb_1
XFILLER_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output444_A _1919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1762__A _1762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1201_ _1221_/A vssd1 vssd1 vccd1 vccd1 _1208_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_output611_A _1743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1512__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1132_ _1132_/A vssd1 vssd1 vccd1 vccd1 _1132_/X sky130_fd_sc_hd__buf_2
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1063_ _1733_/A _2151_/Q _1760_/A vssd1 vssd1 vccd1 vccd1 _1064_/A sky130_fd_sc_hd__and3_1
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2117__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1965_ _1964_/X _1965_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0916_ _1732_/A _1709_/A vssd1 vssd1 vccd1 vccd1 _0917_/A sky130_fd_sc_hd__and2_1
X_1896_ _0888_/X _1896_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1896_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0847_ _2154_/Q vssd1 vssd1 vccd1 vccd1 _1148_/A sky130_fd_sc_hd__inv_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput209 wr_data[124] vssd1 vssd1 vccd1 vccd1 _0997_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1503__B1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_33_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input175_A read_interactive_req_core0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input36_A core0_data_print[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0926__A _0926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output394_A _1701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1750_ _1750_/A vssd1 vssd1 vccd1 vccd1 _1750_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1757__A _1757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1981__A0 _1980_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output561_A _2106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1681_ _1681_/A vssd1 vssd1 vccd1 vccd1 _1681_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1115_ _2019_/Q _1115_/B vssd1 vssd1 vccd1 vccd1 _1116_/A sky130_fd_sc_hd__and2_1
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2095_ _2149_/CLK _2095_/D vssd1 vssd1 vccd1 vccd1 _2095_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1046_ _1046_/A vssd1 vssd1 vccd1 vccd1 _1046_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1948_ _0944_/X _1948_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1948_/X sky130_fd_sc_hd__mux2_2
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1879_ _1878_/X _1336_/A _1954_/S vssd1 vssd1 vccd1 vccd1 _1879_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input292_A wr_data[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1963__A0 _1962_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1487__A _1487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1802_ _1801_/X _1685_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1802_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1954__A0 _1953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1733_ _1733_/A vssd1 vssd1 vccd1 vccd1 _1733_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_113_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2147_ _1767_/X _2147_/D vssd1 vssd1 vccd1 vccd1 _2147_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2078_ _1767_/X _2078_/D vssd1 vssd1 vccd1 vccd1 _2078_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1029_ _1733_/A _2151_/Q _1743_/A vssd1 vssd1 vccd1 vccd1 _1030_/A sky130_fd_sc_hd__and3_1
XFILLER_50_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_22_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input138_A la_data_in[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1476__A2 _1470_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input305_A wr_data[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1400__A2 _1396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1380_ _2121_/Q _1373_/X input78/X _1376_/X vssd1 vssd1 vccd1 vccd1 _2121_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1164__A1 _2152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output524_A _2072_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2001_ _2000_/X _2001_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _2001_/X sky130_fd_sc_hd__mux2_4
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1467__A2 _1438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1716_ _1716_/A vssd1 vssd1 vccd1 vccd1 _1716_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_104_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1155__B2 _1150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1458__A2 _1452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1918__A0 _1917_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1394__A1 _2131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1671__778 vssd1 vssd1 vccd1 vccd1 _1671__778/HI la_data_out[120] sky130_fd_sc_hd__conb_1
XFILLER_123_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input255_A wr_data[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_77_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0918__B _0930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1565__672 vssd1 vssd1 vccd1 vccd1 _1565__672/HI la_data_out[13] sky130_fd_sc_hd__conb_1
XFILLER_14_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0880_ _0880_/A vssd1 vssd1 vccd1 vccd1 _0880_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1765__A _1765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2150__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output474_A _2142_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1385__A1 _2124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1501_ _1508_/A vssd1 vssd1 vccd1 vccd1 _1501_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output641_A _1084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1432_ _1439_/A vssd1 vssd1 vccd1 vccd1 _1432_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1363_ _2113_/Q _1357_/X input72/X _1360_/X vssd1 vssd1 vccd1 vccd1 _2113_/D sky130_fd_sc_hd__a22o_1
X_1294_ _1297_/A _1303_/A _1293_/Y vssd1 vssd1 vccd1 vccd1 _1294_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1005__A _1005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput630 _1122_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_105_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput641 _1084_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XFILLER_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2023__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input66_A dout0_to_sram[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output591_A _1735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ _1980_/X _1981_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1981_/X sky130_fd_sc_hd__mux2_2
X_0932_ _1732_/A _1713_/A vssd1 vssd1 vccd1 vccd1 _0933_/A sky130_fd_sc_hd__and2_1
XFILLER_9_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0863_ _0863_/A vssd1 vssd1 vccd1 vccd1 _2018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1415_ _2146_/Q _1410_/X input73/X _1411_/X vssd1 vssd1 vccd1 vccd1 _2146_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2046__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1346_ _1346_/A _1346_/B vssd1 vssd1 vccd1 vccd1 _1347_/A sky130_fd_sc_hd__or2_1
XFILLER_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1530__A1 _2096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1277_ _1277_/A _1277_/B vssd1 vssd1 vccd1 vccd1 _1289_/B sky130_fd_sc_hd__or2_1
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_137_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput471 _2140_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[118] sky130_fd_sc_hd__buf_2
XFILLER_121_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput460 _2130_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[108] sky130_fd_sc_hd__buf_2
Xoutput482 _2034_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput493 _2044_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1521__A1 _2089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input120_A la_data_in[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input218_A wr_data[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1677__784 vssd1 vssd1 vccd1 vccd1 _1677__784/HI la_data_out[126] sky130_fd_sc_hd__conb_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2069__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1200_ _1204_/A vssd1 vssd1 vccd1 vccd1 _1221_/A sky130_fd_sc_hd__inv_2
XANTENNA__1512__A1 _2082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output604_A _1765_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1131_ _2019_/Q _1131_/B vssd1 vssd1 vccd1 vccd1 _1132_/A sky130_fd_sc_hd__and2_1
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1062_ _1062_/A vssd1 vssd1 vccd1 vccd1 _1062_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1964_ _0961_/X _1964_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1964_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0915_ _0915_/A vssd1 vssd1 vccd1 vccd1 _0915_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1895_ _1894_/X _0882_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1895_/X sky130_fd_sc_hd__mux2_4
X_0846_ _0870_/B _0875_/C vssd1 vssd1 vccd1 vccd1 _2017_/S sky130_fd_sc_hd__nor2_2
XFILLER_127_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1503__A1 _2075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1329_ _1343_/A _1329_/B vssd1 vssd1 vccd1 vccd1 _1341_/B sky130_fd_sc_hd__or2_1
XFILLER_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1990__A1 _1990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input168_A la_data_in[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input29_A core0_data_print[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1802__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0926__B _0930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1605__712 vssd1 vssd1 vccd1 vccd1 _1605__712/HI la_data_out[53] sky130_fd_sc_hd__conb_1
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1103__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1981__A1 _1981_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1430__B1 _2026_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1680_ _1680_/A vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_output554_A _2100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1497__B1 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_54_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1114_ _1114_/A vssd1 vssd1 vccd1 vccd1 _1114_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2094_ _2149_/CLK _2094_/D vssd1 vssd1 vccd1 vccd1 _2094_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1013__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1045_ _1733_/A _2151_/Q _1751_/A vssd1 vssd1 vccd1 vccd1 _1046_/A sky130_fd_sc_hd__and3_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1947_ _1946_/X _0938_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1947_/X sky130_fd_sc_hd__mux2_4
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1972__A1 _1972_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1878_ _1877_/X _1340_/Y _2013_/S vssd1 vssd1 vccd1 vccd1 _1878_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1488__B1 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input285_A wr_data[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1412__B1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2107__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0937__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1801_ _1800_/X _1189_/A _1922_/S vssd1 vssd1 vccd1 vccd1 _1801_/X sky130_fd_sc_hd__mux2_1
X_1732_ _1732_/A vssd1 vssd1 vccd1 vccd1 _1732_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1954__A1 _1954_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0847__A _2154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2146_ _1767_/X _2146_/D vssd1 vssd1 vccd1 vccd1 _2146_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1890__A0 _1889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2077_ _2149_/CLK _2077_/D vssd1 vssd1 vccd1 vccd1 _2077_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1582__689 vssd1 vssd1 vccd1 vccd1 _1582__689/HI la_data_out[30] sky130_fd_sc_hd__conb_1
X_1028_ _1028_/A vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__buf_2
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_18_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input200_A wr_data[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input96_A la_data_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1936__A1 _1936_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1164__A2 _1150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2000_ _0998_/X _2000_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _2000_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1715_ _1715_/A vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2129_ _2149_/CLK _2129_/D vssd1 vssd1 vccd1 vccd1 _2129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_82_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1900__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1918__A1 _1918_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input150_A la_data_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input248_A wr_data[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input11_A addr_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1810__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1111__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1909__A1 _1909_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output467_A _2136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1500_ _1507_/A vssd1 vssd1 vccd1 vccd1 _1500_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1431_ _1438_/A vssd1 vssd1 vccd1 vccd1 _1431_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1362_ _2112_/Q _1357_/X input71/X _1360_/X vssd1 vssd1 vccd1 vccd1 _2112_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1293_ _1297_/A _1303_/A vssd1 vssd1 vccd1 vccd1 _1293_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput190 wr_data[107] vssd1 vssd1 vccd1 vccd1 _0926_/A sky130_fd_sc_hd__buf_2
XANTENNA__1005__B _1009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1021__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput620 _1104_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
Xoutput642 _1086_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput631 _1124_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1691__A _1691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input3_A addr_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1588__695 vssd1 vssd1 vccd1 vccd1 _1588__695/HI la_data_out[36] sky130_fd_sc_hd__conb_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2013__A0 _2012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input198_A wr_data[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input59_A dout0_to_sram[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1805__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_133_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0945__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1980_ _0978_/X _1980_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1980_/X sky130_fd_sc_hd__mux2_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ _0931_/A vssd1 vssd1 vccd1 vccd1 _0931_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_output584_A _1747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0862_ _2016_/X _1139_/B _2019_/Q vssd1 vssd1 vccd1 vccd1 _0863_/A sky130_fd_sc_hd__or3_1
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_115_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1414_ _2145_/Q _1410_/X input72/X _1411_/X vssd1 vssd1 vccd1 vccd1 _2145_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1345_ _1341_/A _1332_/X _1344_/Y vssd1 vssd1 vccd1 vccd1 _1345_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1276_ _1274_/A _1274_/B _1275_/Y vssd1 vssd1 vccd1 vccd1 _1276_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1622__729 vssd1 vssd1 vccd1 vccd1 _1622__729/HI la_data_out[70] sky130_fd_sc_hd__conb_1
XFILLER_12_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1686__A _1686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput461 _2131_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[109] sky130_fd_sc_hd__buf_2
Xoutput450 _2019_/Q vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_2
XFILLER_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput472 _2141_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[119] sky130_fd_sc_hd__buf_2
Xoutput494 _2045_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[23] sky130_fd_sc_hd__buf_2
Xoutput483 _2035_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_120_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2140__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input113_A la_data_in[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_129_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output332_A _1691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1130_ _1130_/A vssd1 vssd1 vccd1 vccd1 _1130_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1061_ _1733_/A _2151_/Q _1759_/A vssd1 vssd1 vccd1 vccd1 _1062_/A sky130_fd_sc_hd__and3_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1963_ _1962_/X _0954_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1963_/X sky130_fd_sc_hd__mux2_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_0914_ _0914_/A _0930_/B vssd1 vssd1 vccd1 vccd1 _0915_/A sky130_fd_sc_hd__and2_1
X_1894_ _1893_/X _1894_/A1 _1990_/S vssd1 vssd1 vccd1 vccd1 _1894_/X sky130_fd_sc_hd__mux2_4
X_0845_ _2155_/Q _0841_/X _2153_/Q _0852_/B vssd1 vssd1 vccd1 vccd1 _2153_/D sky130_fd_sc_hd__o211a_1
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1328_ input9/X _1315_/Y _1338_/B vssd1 vssd1 vccd1 vccd1 _1328_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1259_ input3/X _1248_/Y _1269_/B vssd1 vssd1 vccd1 vccd1 _1259_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_133_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input230_A wr_data[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1644__751 vssd1 vssd1 vccd1 vccd1 _1644__751/HI la_data_out[92] sky130_fd_sc_hd__conb_1
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1103__B _1103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2036__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1430__A1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1430__B2 _1425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output547_A _2093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1497__A1 _2071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2093_ _1767_/X _2093_/D vssd1 vssd1 vccd1 vccd1 _2093_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1113_ _2019_/Q _1113_/B vssd1 vssd1 vccd1 vccd1 _1114_/A sky130_fd_sc_hd__and2_1
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1044_ _1044_/A vssd1 vssd1 vccd1 vccd1 _1044_/X sky130_fd_sc_hd__buf_6
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1013__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1946_ _1945_/X _1946_/A1 _2010_/S vssd1 vssd1 vccd1 vccd1 _1946_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1877_ _1876_/X _1342_/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1877_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1903__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1628__735 vssd1 vssd1 vccd1 vccd1 _1628__735/HI la_data_out[76] sky130_fd_sc_hd__conb_1
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2059__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1412__A1 _2143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input278_A wr_data[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input180_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input41_A core0_data_print[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1813__S _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0937__B _1714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0953__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output497_A _2048_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1800_ _1799_/X _1192_/Y _2013_/S vssd1 vssd1 vccd1 vccd1 _1800_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1731_ _1731_/A vssd1 vssd1 vccd1 vccd1 _1731_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _1767_/X _2145_/D vssd1 vssd1 vccd1 vccd1 _2145_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1890__A1 _1890_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2076_ _1767_/X _2076_/D vssd1 vssd1 vccd1 vccd1 _2076_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1027_ _1733_/A _2151_/Q _1742_/A vssd1 vssd1 vccd1 vccd1 _1028_/A sky130_fd_sc_hd__and3_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1929_ _1928_/X _1929_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1929_/X sky130_fd_sc_hd__mux2_2
XANTENNA__1694__A _1694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input89_A la_data_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1808__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1109__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output412_A _1707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1388__B1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1714_ _1714_/A vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1019__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0858__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_98_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2128_ _2149_/CLK _2128_/D vssd1 vssd1 vccd1 vccd1 _2128_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ _2155_/CLK _2059_/D vssd1 vssd1 vccd1 vccd1 _2059_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1379__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_135_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_131_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input143_A la_data_in[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_122_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1111__B _1111_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output362_A _1014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1430_ input79/X _1422_/X _2026_/Q _1425_/X vssd1 vssd1 vccd1 vccd1 _2026_/D sky130_fd_sc_hd__o22a_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1361_ _2111_/Q _1357_/X input70/X _1360_/X vssd1 vssd1 vccd1 vccd1 _2111_/D sky130_fd_sc_hd__a22o_1
XFILLER_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1542__B1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output627_A _1116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1292_ _1302_/A vssd1 vssd1 vccd1 vccd1 _1297_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput180 wb_rst_i vssd1 vssd1 vccd1 vccd1 _2016_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput191 wr_data[108] vssd1 vssd1 vccd1 vccd1 _0930_/A sky130_fd_sc_hd__buf_2
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1021__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput610 _1742_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[8] sky130_fd_sc_hd__buf_2
Xoutput621 _1106_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput632 _1126_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput643 _1088_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1911__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_136_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2013__A1 _2013_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input260_A wr_data[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1524__B1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1821__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0945__B _1716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_45_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0930_ _0930_/A _0930_/B vssd1 vssd1 vccd1 vccd1 _0931_/A sky130_fd_sc_hd__and2_2
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output577_A _2121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0861_ _0861_/A vssd1 vssd1 vccd1 vccd1 _1139_/B sky130_fd_sc_hd__inv_2
XFILLER_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1515__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1413_ _2144_/Q _1410_/X input71/X _1411_/X vssd1 vssd1 vccd1 vccd1 _2144_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1344_ _1344_/A vssd1 vssd1 vccd1 vccd1 _1344_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_84_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1275_ _1319_/D vssd1 vssd1 vccd1 vccd1 _1275_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1661__768 vssd1 vssd1 vccd1 vccd1 _1661__768/HI la_data_out[110] sky130_fd_sc_hd__conb_1
XFILLER_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0871__A _2154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2092__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1555__662 vssd1 vssd1 vccd1 vccd1 _1555__662/HI la_data_out[3] sky130_fd_sc_hd__conb_1
XANTENNA__1906__S _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput462 _2032_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[10] sky130_fd_sc_hd__buf_2
Xoutput451 _2022_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[0] sky130_fd_sc_hd__buf_2
Xoutput440 _1903_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[3] sky130_fd_sc_hd__buf_2
Xoutput495 _2046_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[24] sky130_fd_sc_hd__buf_2
Xoutput473 _2033_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1506__B1 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput484 _2036_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input106_A la_data_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1993__A0 _1992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input71_A dout0_to_sram[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1816__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1117__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0956__A _0956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output325_A _1803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1060_ _1060_/A vssd1 vssd1 vccd1 vccd1 _1060_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1962_ _1961_/X _1962_/A1 _1990_/S vssd1 vssd1 vccd1 vccd1 _1962_/X sky130_fd_sc_hd__mux2_4
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0913_ _0976_/A vssd1 vssd1 vccd1 vccd1 _0930_/B sky130_fd_sc_hd__buf_2
X_1893_ _1892_/X _1893_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1893_/X sky130_fd_sc_hd__mux2_1
X_0844_ _0841_/X _0875_/C _0866_/A _2017_/X _0852_/B vssd1 vssd1 vccd1 vccd1 _2154_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1027__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1327_ _1343_/A _1327_/B vssd1 vssd1 vccd1 vccd1 _1338_/B sky130_fd_sc_hd__or2_1
XFILLER_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1258_ _1263_/A _1265_/A _1258_/C vssd1 vssd1 vccd1 vccd1 _1269_/B sky130_fd_sc_hd__or3_1
X_1189_ _1189_/A vssd1 vssd1 vccd1 vccd1 _1212_/B sky130_fd_sc_hd__inv_2
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1697__A _1697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1975__A0 _1974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA_input223_A wr_data[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1430__A2 _1422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2092_ _2149_/CLK _2092_/D vssd1 vssd1 vccd1 vccd1 _2092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1112_ _1112_/A vssd1 vssd1 vccd1 vccd1 _1112_/X sky130_fd_sc_hd__clkbuf_2
X_1043_ _1733_/A _2151_/Q _1750_/A vssd1 vssd1 vccd1 vccd1 _1044_/A sky130_fd_sc_hd__and3_1
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1013__C _1735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1945_ _1944_/X _1945_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1945_/X sky130_fd_sc_hd__mux2_2
XFILLER_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1957__A0 _1956_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1876_ _1336_/A _1345_/Y _1882_/S vssd1 vssd1 vccd1 vccd1 _1876_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2130__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1185__A1 _1177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1667__774 vssd1 vssd1 vccd1 vccd1 _1667__774/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_119_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input173_A la_oenb[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input34_A core0_data_print[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output392_A _1718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2153__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1730_ _1730_/A vssd1 vssd1 vccd1 vccd1 _1730_/X sky130_fd_sc_hd__buf_2
XFILLER_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_131_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _1767_/X _2144_/D vssd1 vssd1 vccd1 vccd1 _2144_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_39_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2075_ _1767_/X _2075_/D vssd1 vssd1 vccd1 vccd1 _2075_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1026_ _1026_/A vssd1 vssd1 vccd1 vccd1 _1026_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1928_ _0923_/X _1928_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1928_/X sky130_fd_sc_hd__mux2_8
XFILLER_135_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1859_ _1858_/X _1307_/Y _2012_/S vssd1 vssd1 vccd1 vccd1 _1859_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1914__S _1934_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2021__D _2152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2026__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input290_A wr_data[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_113_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1109__B _1109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1824__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1125__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1388__A1 _2127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1713_ _1713_/A vssd1 vssd1 vccd1 vccd1 _1713_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_132_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1019__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2049__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0858__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1035__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2127_ _1767_/X _2127_/D vssd1 vssd1 vccd1 vccd1 _2127_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2155_/CLK _2058_/D vssd1 vssd1 vccd1 vccd1 _2058_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1009_ _1009_/A _1009_/B vssd1 vssd1 vccd1 vccd1 _1010_/A sky130_fd_sc_hd__and2_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1909__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_6_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1379__A1 _2120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input136_A la_data_in[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input303_A wr_data[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1819__S _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1572__679 vssd1 vssd1 vccd1 vccd1 _1572__679/HI la_data_out[20] sky130_fd_sc_hd__conb_1
X_1360_ _1520_/A vssd1 vssd1 vccd1 vccd1 _1360_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1542__A1 _2104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output522_A _2071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1291_ input6/X vssd1 vssd1 vccd1 vccd1 _1302_/A sky130_fd_sc_hd__inv_2
Xinput170 la_data_in[98] vssd1 vssd1 vccd1 vccd1 _1732_/A sky130_fd_sc_hd__buf_12
XFILLER_76_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput181 we vssd1 vssd1 vccd1 vccd1 _1146_/B sky130_fd_sc_hd__clkbuf_1
Xinput192 wr_data[109] vssd1 vssd1 vccd1 vccd1 _0935_/A sky130_fd_sc_hd__buf_2
XFILLER_64_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1021__C _1739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_117_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput600 _1762_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[28] sky130_fd_sc_hd__buf_2
Xoutput611 _1743_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[9] sky130_fd_sc_hd__buf_2
Xoutput644 _1090_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput633 _1128_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
Xoutput622 _1108_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
XFILLER_99_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1489_ _2065_/Q _1486_/X input55/X _1487_/X vssd1 vssd1 vccd1 vccd1 _2065_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_52_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input253_A wr_data[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1524__A1 _2092_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0860_ _0857_/Y _2150_/Q _2016_/X _0859_/X vssd1 vssd1 vccd1 vccd1 _2150_/D sky130_fd_sc_hd__a211o_1
XANTENNA_output472_A _2141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1412_ _2143_/Q _1410_/X input70/X _1411_/X vssd1 vssd1 vccd1 vccd1 _2143_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1515__B2 _1487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1515__A1 _2085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1343_ _1343_/A _1346_/A _1343_/C vssd1 vssd1 vccd1 vccd1 _1344_/A sky130_fd_sc_hd__or3_1
XFILLER_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1274_ _1274_/A _1274_/B vssd1 vssd1 vccd1 vccd1 _1319_/D sky130_fd_sc_hd__or2_1
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0871__B _2152_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1451__B1 _2041_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0989_ _0989_/A _0993_/B vssd1 vssd1 vccd1 vccd1 _0990_/A sky130_fd_sc_hd__and2_1
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
Xoutput452 _2122_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[100] sky130_fd_sc_hd__buf_2
XFILLER_133_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput430 _1983_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[23] sky130_fd_sc_hd__buf_2
Xoutput441 _1907_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[4] sky130_fd_sc_hd__buf_2
Xoutput463 _2132_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[110] sky130_fd_sc_hd__buf_2
XANTENNA__1506__A1 _2078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput496 _2047_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[25] sky130_fd_sc_hd__buf_2
Xoutput485 _2037_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[15] sky130_fd_sc_hd__buf_2
Xoutput474 _2142_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[120] sky130_fd_sc_hd__buf_2
XFILLER_120_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1922__S _1922_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1223__A _1223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1442__B1 _2034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1993__A1 _1993_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input64_A dout0_to_sram[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1117__B _1117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1832__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0956__B _0972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1133__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output318_A _1875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0972__A _0972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ _1960_/X _1961_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1961_/X sky130_fd_sc_hd__mux2_1
X_1892_ _0884_/X _1892_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1892_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0912_ _0912_/A vssd1 vssd1 vccd1 vccd1 _0912_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1433__B1 _2027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1578__685 vssd1 vssd1 vccd1 vccd1 _1578__685/HI la_data_out[26] sky130_fd_sc_hd__conb_1
X_0843_ _2016_/X _0843_/B vssd1 vssd1 vccd1 vccd1 _0852_/B sky130_fd_sc_hd__nor2_2
XFILLER_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_102_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1027__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1326_ _1334_/A vssd1 vssd1 vccd1 vccd1 _1343_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1043__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1257_ input3/X vssd1 vssd1 vccd1 vccd1 _1265_/A sky130_fd_sc_hd__inv_2
X_1188_ _1212_/A _1186_/B _1187_/Y vssd1 vssd1 vccd1 vccd1 _1188_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1917__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input216_A wr_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_90_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1415__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1966__A1 _1966_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1827__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1612__719 vssd1 vssd1 vccd1 vccd1 _1612__719/HI la_data_out[60] sky130_fd_sc_hd__conb_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2082__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output435_A _2003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2091_ _1767_/X _2091_/D vssd1 vssd1 vccd1 vccd1 _2091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1111_ _2019_/Q _1111_/B vssd1 vssd1 vccd1 vccd1 _1112_/A sky130_fd_sc_hd__and2_1
XFILLER_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1042_ _1042_/A vssd1 vssd1 vccd1 vccd1 _1042_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1406__B1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1944_ _0940_/X _1944_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1944_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1875_ _1335_/X _1874_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1875_/X sky130_fd_sc_hd__mux2_4
XFILLER_116_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0877__A _0891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1309_ input7/X _1297_/Y _1308_/X vssd1 vssd1 vccd1 vccd1 _1309_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1948__A1 _1948_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input166_A la_data_in[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input27_A core0_data_print[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_16_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output385_A _1711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output552_A _2098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _1767_/X _2143_/D vssd1 vssd1 vccd1 vccd1 _2143_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2074_ _2155_/CLK _2074_/D vssd1 vssd1 vccd1 vccd1 _2074_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1025_ _1733_/A _2151_/Q _1741_/A vssd1 vssd1 vccd1 vccd1 _1026_/A sky130_fd_sc_hd__and3_1
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1593__700 vssd1 vssd1 vccd1 vccd1 _1593__700/HI la_data_out[41] sky130_fd_sc_hd__conb_1
X_1927_ _1926_/X _0917_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1927_/X sky130_fd_sc_hd__mux2_4
X_1858_ input7/X _1309_/X _1882_/S vssd1 vssd1 vccd1 vccd1 _1858_/X sky130_fd_sc_hd__mux2_1
X_1634__741 vssd1 vssd1 vccd1 vccd1 _1634__741/HI la_data_out[82] sky130_fd_sc_hd__conb_1
X_1789_ _1788_/X _1168_/B _1922_/S vssd1 vssd1 vccd1 vccd1 _1789_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1930__S _1938_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input283_A wr_data[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2001__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1125__B _1125_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1840__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0964__B _0972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2120__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1141__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1618__725 vssd1 vssd1 vccd1 vccd1 _1618__725/HI la_data_out[66] sky130_fd_sc_hd__conb_1
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1712_ _1712_/A vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1019__C _1738_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1035__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2126_ _2149_/CLK _2126_/D vssd1 vssd1 vccd1 vccd1 _2126_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1051__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2155_/CLK _2057_/D vssd1 vssd1 vccd1 vccd1 _2057_/Q sky130_fd_sc_hd__dfxtp_1
X_1008_ _1008_/A vssd1 vssd1 vccd1 vccd1 _1008_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1925__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2143__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_73_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input129_A la_data_in[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input94_A la_data_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2016__A0 _1766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_127_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1835__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_110_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1290_ input5/X _1278_/Y _1310_/A vssd1 vssd1 vccd1 vccd1 _1290_/X sky130_fd_sc_hd__o21a_1
Xinput171 la_data_in[99] vssd1 vssd1 vccd1 vccd1 _1733_/A sky130_fd_sc_hd__buf_12
Xinput160 la_data_in[89] vssd1 vssd1 vccd1 vccd1 _1759_/A sky130_fd_sc_hd__buf_4
XFILLER_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xinput193 wr_data[10] vssd1 vssd1 vccd1 vccd1 _1930_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput182 wr_data[0] vssd1 vssd1 vccd1 vccd1 _1890_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
Xoutput601 _1763_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[29] sky130_fd_sc_hd__buf_2
XFILLER_133_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput623 _1110_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput612 _2017_/S vssd1 vssd1 vccd1 vccd1 ready sky130_fd_sc_hd__buf_2
Xoutput634 _1130_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput645 _1092_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_101_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1488_ _2064_/Q _1486_/X input54/X _1487_/X vssd1 vssd1 vccd1 vccd1 _2064_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0885__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2109_ _2149_/CLK _2109_/D vssd1 vssd1 vccd1 vccd1 _2109_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_117_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input246_A wr_data[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1288__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2039__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output465_A _2134_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1411_ _1411_/A vssd1 vssd1 vccd1 vccd1 _1411_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output632_A _1126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1342_ _1336_/A _1330_/Y _1341_/X vssd1 vssd1 vccd1 vccd1 _1342_/X sky130_fd_sc_hd__o21a_1
XFILLER_95_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1273_ input4/X _1261_/Y _1284_/B vssd1 vssd1 vccd1 vccd1 _1273_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1451__A1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0988_ _0988_/A vssd1 vssd1 vccd1 vccd1 _0988_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput420 _1947_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[14] sky130_fd_sc_hd__buf_2
XFILLER_133_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput453 _2123_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[101] sky130_fd_sc_hd__buf_2
Xoutput431 _1987_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[24] sky130_fd_sc_hd__buf_2
Xoutput442 _1911_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[5] sky130_fd_sc_hd__buf_2
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput475 _2143_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[121] sky130_fd_sc_hd__buf_2
Xoutput464 _2133_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[111] sky130_fd_sc_hd__buf_2
Xoutput486 _2038_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[16] sky130_fd_sc_hd__buf_2
Xoutput497 _2048_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A addr_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1442__A1 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input196_A wr_data[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_10_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_136_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input57_A dout0_to_sram[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1133__B _1133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0972__B _0972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1960_ _0957_/X _1960_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1960_/X sky130_fd_sc_hd__mux2_1
X_1891_ _1890_/X _0865_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1891_/X sky130_fd_sc_hd__mux2_2
X_0911_ _1732_/A _1708_/A vssd1 vssd1 vccd1 vccd1 _0912_/A sky130_fd_sc_hd__and2_1
XANTENNA__1433__A1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_0842_ _2155_/Q _2153_/Q vssd1 vssd1 vccd1 vccd1 _0875_/C sky130_fd_sc_hd__or2_2
XFILLER_115_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1027__C _1742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1325_ input9/X vssd1 vssd1 vccd1 vccd1 _1334_/A sky130_fd_sc_hd__inv_2
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1043__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1256_ _1252_/A _1254_/B _1255_/Y vssd1 vssd1 vccd1 vccd1 _1256_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1187_ _1198_/B vssd1 vssd1 vccd1 vccd1 _1187_/Y sky130_fd_sc_hd__inv_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1933__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input209_A wr_data[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input111_A la_data_in[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1415__A1 _2146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2004__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1651__758 vssd1 vssd1 vccd1 vccd1 _1651__758/HI la_data_out[99] sky130_fd_sc_hd__conb_1
XFILLER_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1843__S _1942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1110_ _1110_/A vssd1 vssd1 vccd1 vccd1 _1110_/X sky130_fd_sc_hd__buf_2
XANTENNA_output428_A _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1351__B1 _1349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2090_ _2149_/CLK _2090_/D vssd1 vssd1 vccd1 vccd1 _2090_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0983__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1041_ _1733_/A _2151_/Q _1749_/A vssd1 vssd1 vccd1 vccd1 _1042_/A sky130_fd_sc_hd__and3_1
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1406__A1 _2139_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1943_ _1942_/X _0933_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1943_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1874_ _1873_/X _1697_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1874_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_115_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_1308_ _1308_/A _1319_/B vssd1 vssd1 vccd1 vccd1 _1308_/X sky130_fd_sc_hd__or2_1
X_1239_ _1239_/A _1239_/B vssd1 vssd1 vccd1 vccd1 _1250_/B sky130_fd_sc_hd__or2_1
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1928__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_121_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input159_A la_data_in[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1838__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_124_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _1767_/X _2142_/D vssd1 vssd1 vccd1 vccd1 _2142_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2073_ _1767_/X _2073_/D vssd1 vssd1 vccd1 vccd1 _2073_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1024_ _1024_/A vssd1 vssd1 vccd1 vccd1 _1024_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1926_ _1925_/X _1926_/A1 _1958_/S vssd1 vssd1 vccd1 vccd1 _1926_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1049__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1857_ _1300_/Y _1856_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1857_/X sky130_fd_sc_hd__mux2_1
X_1673__780 vssd1 vssd1 vccd1 vccd1 _1673__780/HI la_data_out[122] sky130_fd_sc_hd__conb_1
X_1788_ _1787_/X _1169_/Y _2013_/S vssd1 vssd1 vccd1 vccd1 _1788_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_72_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__2072__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_138_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input276_A wr_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1422__A _1438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output495_A _2046_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1657__764 vssd1 vssd1 vccd1 vccd1 _1657__764/HI la_data_out[106] sky130_fd_sc_hd__conb_1
X_1711_ _1711_/A vssd1 vssd1 vccd1 vccd1 _1711_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1545__B1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1035__C _1746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2125_ _2149_/CLK _2125_/D vssd1 vssd1 vccd1 vccd1 _2125_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_54_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2056_ _2155_/CLK _2056_/D vssd1 vssd1 vccd1 vccd1 _2056_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1007_ _1732_/A _1731_/A vssd1 vssd1 vccd1 vccd1 _1008_/A sky130_fd_sc_hd__and2_1
XANTENNA__1051__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2095__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1909_ _1908_/X _1909_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1909_/X sky130_fd_sc_hd__mux2_4
XFILLER_135_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1536__B1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1941__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input87_A la_data_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2012__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1851__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput161 la_data_in[8] vssd1 vssd1 vccd1 vccd1 _1688_/A sky130_fd_sc_hd__buf_4
Xinput150 la_data_in[7] vssd1 vssd1 vccd1 vccd1 _1687_/A sky130_fd_sc_hd__buf_4
XFILLER_95_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput172 la_data_in[9] vssd1 vssd1 vccd1 vccd1 _1689_/A sky130_fd_sc_hd__clkbuf_2
Xinput194 wr_data[110] vssd1 vssd1 vccd1 vccd1 _0939_/A sky130_fd_sc_hd__clkbuf_1
Xinput183 wr_data[100] vssd1 vssd1 vccd1 vccd1 _0897_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0991__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput602 _1736_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[2] sky130_fd_sc_hd__buf_2
XFILLER_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1518__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput624 _1112_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput613 _1766_/X vssd1 vssd1 vccd1 vccd1 reset_core sky130_fd_sc_hd__buf_2
Xoutput635 _1132_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
Xoutput646 _1094_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1487_ _1487_/A vssd1 vssd1 vccd1 vccd1 _1487_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0885__B _1702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ _2149_/CLK _2108_/D vssd1 vssd1 vccd1 vccd1 _2108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2039_ _2155_/CLK _2039_/D vssd1 vssd1 vccd1 vccd1 _2039_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1936__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2110__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1509__B1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input239_A wr_data[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input141_A la_data_in[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_100_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1700__A _1700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2007__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1846__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1410_ _1410_/A vssd1 vssd1 vccd1 vccd1 _1410_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output625_A _1114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1341_ _1341_/A _1341_/B vssd1 vssd1 vccd1 vccd1 _1341_/X sky130_fd_sc_hd__or2_1
XFILLER_95_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1272_ _1277_/A _1272_/B vssd1 vssd1 vccd1 vccd1 _1284_/B sky130_fd_sc_hd__or2_1
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1987__A0 _1986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0987_ _1732_/A _1726_/A vssd1 vssd1 vccd1 vccd1 _0988_/A sky130_fd_sc_hd__and2_1
XANTENNA__2133__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput410 _1705_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[5] sky130_fd_sc_hd__buf_2
Xoutput443 _1915_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[6] sky130_fd_sc_hd__buf_2
XFILLER_133_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput432 _1991_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[25] sky130_fd_sc_hd__buf_2
XANTENNA__1057__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput421 _1951_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[15] sky130_fd_sc_hd__buf_2
Xoutput476 _2144_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[122] sky130_fd_sc_hd__buf_2
Xoutput454 _2124_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[102] sky130_fd_sc_hd__buf_2
Xoutput465 _2134_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[112] sky130_fd_sc_hd__buf_2
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput487 _2039_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[17] sky130_fd_sc_hd__buf_2
X_1539_ _2103_/Q _1533_/X input61/X _1534_/X vssd1 vssd1 vccd1 vccd1 _2103_/D sky130_fd_sc_hd__a22o_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput498 _2049_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
X_1562__669 vssd1 vssd1 vccd1 vccd1 _1562__669/HI la_data_out[10] sky130_fd_sc_hd__conb_1
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input189_A wr_data[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1902__A0 _1901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0910_ _0910_/A vssd1 vssd1 vccd1 vccd1 _0910_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1969__A0 _1968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1890_ _1889_/X _1890_/A1 _1934_/S vssd1 vssd1 vccd1 vccd1 _1890_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output575_A _2119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0841_ _0870_/B vssd1 vssd1 vccd1 vccd1 _0841_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1324_ _1319_/C _1322_/B _1323_/Y vssd1 vssd1 vccd1 vccd1 _1324_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1255_ _1265_/B vssd1 vssd1 vccd1 vccd1 _1255_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1043__C _1750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1186_ _1186_/A _1186_/B vssd1 vssd1 vccd1 vccd1 _1198_/B sky130_fd_sc_hd__or2_1
XFILLER_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_80_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_118_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2029__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_75_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_130_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input104_A la_data_in[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_137_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1425__A _1439_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1351__A1 _1336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0983__B _1725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1040_ _1040_/A vssd1 vssd1 vccd1 vccd1 _1040_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1584__691 vssd1 vssd1 vccd1 vccd1 _1584__691/HI la_data_out[32] sky130_fd_sc_hd__conb_1
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1942_ _1941_/X _1942_/A1 _1942_/S vssd1 vssd1 vccd1 vccd1 _1942_/X sky130_fd_sc_hd__mux2_1
X_1873_ _1872_/X input9/X _1954_/S vssd1 vssd1 vccd1 vccd1 _1873_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_116_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1342__A1 _1336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1307_ _1305_/A _1305_/B _1306_/Y vssd1 vssd1 vccd1 vccd1 _1307_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__0893__B _0909_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1238_ _1235_/A _1226_/Y _1258_/C vssd1 vssd1 vccd1 vccd1 _1238_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1169_ _1175_/B _1157_/Y _1179_/A vssd1 vssd1 vccd1 vccd1 _1169_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_114_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1944__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_69_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1333__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1568__675 vssd1 vssd1 vccd1 vccd1 _1568__675/HI la_data_out[16] sky130_fd_sc_hd__conb_1
XANTENNA_input221_A wr_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2015__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1854__S _2013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_113_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output440_A _1903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output538_A _2085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0994__A _0994_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2141_ _2149_/CLK _2141_/D vssd1 vssd1 vccd1 vccd1 _2141_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2072_ _1767_/X _2072_/D vssd1 vssd1 vccd1 vccd1 _2072_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1023_ _1733_/A _2151_/Q _1740_/A vssd1 vssd1 vccd1 vccd1 _1024_/A sky130_fd_sc_hd__and3_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1925_ _1924_/X _1925_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1925_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1856_ _1855_/X _1694_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1856_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1049__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1787_ _1786_/X _1171_/Y _2012_/S vssd1 vssd1 vccd1 vccd1 _1787_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1065__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1602__709 vssd1 vssd1 vccd1 vccd1 _1602__709/HI la_data_out[50] sky130_fd_sc_hd__conb_1
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_41_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1939__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input171_A la_data_in[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input269_A wr_data[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input32_A core0_data_print[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1703__A _1703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1490__B1 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1849__S _1942_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output488_A _2040_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output390_A _1716_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1710_ _1710_/A vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1545__A1 _2107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _2149_/CLK _2124_/D vssd1 vssd1 vccd1 vccd1 _2124_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_26_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2055_ _2155_/CLK _2055_/D vssd1 vssd1 vccd1 vccd1 _2055_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1006_ _1006_/A vssd1 vssd1 vccd1 vccd1 _1006_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1051__C _1754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1481__B1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1908_ _0902_/X _1908_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1908_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__0899__A _1732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1839_ _1266_/X _1838_/X _1887_/S vssd1 vssd1 vccd1 vccd1 _1839_/X sky130_fd_sc_hd__mux2_4
XFILLER_135_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1536__B2 _1534_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1536__A1 _2100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_1_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput162 la_data_in[90] vssd1 vssd1 vccd1 vccd1 _1760_/A sky130_fd_sc_hd__buf_2
Xinput151 la_data_in[80] vssd1 vssd1 vccd1 vccd1 _1750_/A sky130_fd_sc_hd__clkbuf_2
Xinput140 la_data_in[70] vssd1 vssd1 vccd1 vccd1 _1740_/A sky130_fd_sc_hd__buf_4
Xinput173 la_oenb[96] vssd1 vssd1 vccd1 vccd1 _1767_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xinput195 wr_data[111] vssd1 vssd1 vccd1 vccd1 _0943_/A sky130_fd_sc_hd__buf_2
Xinput184 wr_data[101] vssd1 vssd1 vccd1 vccd1 _0901_/A sky130_fd_sc_hd__buf_2
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output403_A _1728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0991__B _1727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1624__731 vssd1 vssd1 vccd1 vccd1 _1624__731/HI la_data_out[72] sky130_fd_sc_hd__conb_1
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1463__B1 _2049_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput636 _1134_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XANTENNA__1518__A1 _2088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput603 _1764_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[30] sky130_fd_sc_hd__buf_2
Xoutput625 _1114_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput614 _2016_/X vssd1 vssd1 vccd1 vccd1 rst sky130_fd_sc_hd__buf_2
XFILLER_132_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput647 _1768_/X vssd1 vssd1 vccd1 vccd1 we_to_sram sky130_fd_sc_hd__buf_2
XFILLER_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1486_ _1486_/A vssd1 vssd1 vccd1 vccd1 _1486_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2062__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
X_2107_ _2149_/CLK _2107_/D vssd1 vssd1 vccd1 vccd1 _2107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _2155_/CLK _2038_/D vssd1 vssd1 vccd1 vccd1 _2038_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1454__B1 _2042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XANTENNA__1509__A1 _2079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1952__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input134_A la_data_in[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1608__715 vssd1 vssd1 vccd1 vccd1 _1608__715/HI la_data_out[56] sky130_fd_sc_hd__conb_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input301_A wr_data[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2085__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1862__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1340_ _1341_/A _1338_/B _1339_/Y vssd1 vssd1 vccd1 vccd1 _1340_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_96_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1920__A1 _1920_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output520_A _2069_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output618_A _1100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1271_ _1274_/A _1269_/B _1270_/Y vssd1 vssd1 vccd1 vccd1 _1271_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0986_ _0986_/A vssd1 vssd1 vccd1 vccd1 _0986_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput411 _1706_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[6] sky130_fd_sc_hd__buf_2
Xoutput400 _1725_/X vssd1 vssd1 vccd1 vccd1 data_to_core_mem[25] sky130_fd_sc_hd__buf_2
Xoutput433 _1995_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[26] sky130_fd_sc_hd__buf_2
XFILLER_133_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1057__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput422 _1955_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[16] sky130_fd_sc_hd__buf_2
Xoutput444 _1919_/X vssd1 vssd1 vccd1 vccd1 din0_to_sram[7] sky130_fd_sc_hd__buf_2
Xoutput477 _2145_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[123] sky130_fd_sc_hd__buf_2
Xoutput455 _2125_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[103] sky130_fd_sc_hd__buf_2
Xoutput466 _2135_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[113] sky130_fd_sc_hd__buf_2
XANTENNA__1772__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1538_ _2102_/Q _1533_/X input60/X _1534_/X vssd1 vssd1 vccd1 vccd1 _2102_/D sky130_fd_sc_hd__a22o_1
Xoutput488 _2040_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[18] sky130_fd_sc_hd__buf_2
Xoutput499 _2050_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[28] sky130_fd_sc_hd__buf_2
X_1469_ _1507_/A vssd1 vssd1 vccd1 vccd1 _1486_/A sky130_fd_sc_hd__buf_2
XFILLER_87_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1073__A _1733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1978__A1 _1978_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1947__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input251_A wr_data[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1902__A1 _1902_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1711__A _1711_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1418__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1857__S _1887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0840_ _2154_/Q _2152_/Q vssd1 vssd1 vccd1 vccd1 _0870_/B sky130_fd_sc_hd__or2_2
XANTENNA_output470_A _2139_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output568_A _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0997__A _0997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1323_ _1334_/B vssd1 vssd1 vccd1 vccd1 _1323_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1254_ _1263_/A _1254_/B vssd1 vssd1 vccd1 vccd1 _1265_/B sky130_fd_sc_hd__or2_1
XFILLER_77_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1185_ _1177_/A _1173_/A _1195_/B vssd1 vssd1 vccd1 vccd1 _1185_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2100__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1409__B1 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_0969_ _0969_/A vssd1 vssd1 vccd1 vccd1 _0969_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input299_A wr_data[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_23_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_99_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input62_A dout0_to_sram[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1706__A _1706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2123__CLK _2149_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_59_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output316_A _1863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1941_ _1940_/X _1941_/A1 _2013_/S vssd1 vssd1 vccd1 vccd1 _1941_/X sky130_fd_sc_hd__mux2_8
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1872_ _1871_/X _1328_/X _2013_/S vssd1 vssd1 vccd1 vccd1 _1872_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1306_ _1317_/B vssd1 vssd1 vccd1 vccd1 _1306_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1237_ _1244_/A _1237_/B vssd1 vssd1 vccd1 vccd1 _1258_/C sky130_fd_sc_hd__or2_1
XFILLER_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1168_ _1168_/A _1168_/B _1168_/C vssd1 vssd1 vccd1 vccd1 _1179_/A sky130_fd_sc_hd__and3_1
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1099_ _2019_/Q _1099_/B vssd1 vssd1 vccd1 vccd1 _1100_/A sky130_fd_sc_hd__and2_1
XFILLER_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2146__CLK _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1960__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_input214_A wr_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_12_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_112_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output433_A _1995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1870__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2140_ _2149_/CLK _2140_/D vssd1 vssd1 vccd1 vccd1 _2140_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_78_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2071_ _2149_/CLK _2071_/D vssd1 vssd1 vccd1 vccd1 _2071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1022_ _1022_/A vssd1 vssd1 vccd1 vccd1 _1022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1924_ _0919_/X _1924_/A1 _2012_/S vssd1 vssd1 vccd1 vccd1 _1924_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2019__CLK _2155_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1855_ _1854_/X input6/X _1942_/S vssd1 vssd1 vccd1 vccd1 _1855_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1049__C _1753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1786_ _1168_/B _1174_/X _1882_/S vssd1 vssd1 vccd1 vccd1 _1786_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA__1065__B _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1780__S _1882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1081__A _2019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1641__748 vssd1 vssd1 vccd1 vccd1 _1641__748/HI la_data_out[89] sky130_fd_sc_hd__conb_1
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_111_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1251__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1955__S _2015_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_20_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input164_A la_data_in[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput300 wr_data[91] vssd1 vssd1 vccd1 vccd1 _1996_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_121_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input25_A core0_data_print[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_129_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1865__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0989__B _0993_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XANTENNA_output550_A _2096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2123_ _2149_/CLK _2123_/D vssd1 vssd1 vccd1 vccd1 _2123_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_4
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2054_ _2155_/CLK _2054_/D vssd1 vssd1 vccd1 vccd1 _2054_/Q sky130_fd_sc_hd__dfxtp_1
X_1005_ _1005_/A _1009_/B vssd1 vssd1 vccd1 vccd1 _1006_/A sky130_fd_sc_hd__and2_2
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1481__A1 _2059_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1775__S _2012_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1907_ _1906_/X _0896_/X _2015_/S vssd1 vssd1 vccd1 vccd1 _1907_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0899__B _1705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1838_ _1837_/X _1691_/A _2015_/S vssd1 vssd1 vccd1 vccd1 _1838_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1536__A2 _1533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1769_ _1145_/X input1/X _2012_/S vssd1 vssd1 vccd1 vccd1 _1769_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input281_A wr_data[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1714__A _1714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput141 la_data_in[71] vssd1 vssd1 vccd1 vccd1 _1741_/A sky130_fd_sc_hd__buf_4
Xinput152 la_data_in[81] vssd1 vssd1 vccd1 vccd1 _1751_/A sky130_fd_sc_hd__buf_2
Xinput130 la_data_in[61] vssd1 vssd1 vccd1 vccd1 _1729_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput163 la_data_in[91] vssd1 vssd1 vccd1 vccd1 _1761_/A sky130_fd_sc_hd__buf_2
Xinput196 wr_data[112] vssd1 vssd1 vccd1 vccd1 _0947_/A sky130_fd_sc_hd__clkbuf_1
Xinput185 wr_data[102] vssd1 vssd1 vccd1 vccd1 _0905_/A sky130_fd_sc_hd__buf_2
XFILLER_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput174 la_oenb[97] vssd1 vssd1 vccd1 vccd1 _2016_/S sky130_fd_sc_hd__buf_4
XFILLER_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1663__770 vssd1 vssd1 vccd1 vccd1 _1663__770/HI la_data_out[112] sky130_fd_sc_hd__conb_1
XANTENNA__1463__A1 input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output598_A _1760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_8
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput604 _1765_/X vssd1 vssd1 vccd1 vccd1 read_value_to_Elpis[31] sky130_fd_sc_hd__buf_2
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput615 _1076_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
Xoutput626 _1078_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput637 _1080_/X vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1485_ _2063_/Q _1479_/X input84/X _1480_/X vssd1 vssd1 vccd1 vccd1 _2063_/D sky130_fd_sc_hd__a22o_1
XFILLER_101_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
.ends

