VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_controller
  CLASS BLOCK ;
  FOREIGN chip_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN addr0_to_sram[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 396.000 0.830 400.000 ;
    END
  END addr0_to_sram[0]
  PIN addr0_to_sram[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 72.120 400.000 72.720 ;
    END
  END addr0_to_sram[10]
  PIN addr0_to_sram[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 396.000 62.470 400.000 ;
    END
  END addr0_to_sram[11]
  PIN addr0_to_sram[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END addr0_to_sram[12]
  PIN addr0_to_sram[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END addr0_to_sram[13]
  PIN addr0_to_sram[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END addr0_to_sram[14]
  PIN addr0_to_sram[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 105.440 400.000 106.040 ;
    END
  END addr0_to_sram[15]
  PIN addr0_to_sram[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END addr0_to_sram[16]
  PIN addr0_to_sram[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 127.200 400.000 127.800 ;
    END
  END addr0_to_sram[17]
  PIN addr0_to_sram[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 133.320 400.000 133.920 ;
    END
  END addr0_to_sram[18]
  PIN addr0_to_sram[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END addr0_to_sram[19]
  PIN addr0_to_sram[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 9.560 400.000 10.160 ;
    END
  END addr0_to_sram[1]
  PIN addr0_to_sram[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END addr0_to_sram[2]
  PIN addr0_to_sram[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END addr0_to_sram[3]
  PIN addr0_to_sram[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 20.440 400.000 21.040 ;
    END
  END addr0_to_sram[4]
  PIN addr0_to_sram[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 396.000 28.890 400.000 ;
    END
  END addr0_to_sram[5]
  PIN addr0_to_sram[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END addr0_to_sram[6]
  PIN addr0_to_sram[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 396.000 44.070 400.000 ;
    END
  END addr0_to_sram[7]
  PIN addr0_to_sram[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END addr0_to_sram[8]
  PIN addr0_to_sram[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 61.240 400.000 61.840 ;
    END
  END addr0_to_sram[9]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END addr_in[0]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 77.560 400.000 78.160 ;
    END
  END addr_in[11]
  PIN addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 396.000 75.810 400.000 ;
    END
  END addr_in[12]
  PIN addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 85.040 400.000 85.640 ;
    END
  END addr_in[13]
  PIN addr_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.920 400.000 96.520 ;
    END
  END addr_in[14]
  PIN addr_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 107.480 400.000 108.080 ;
    END
  END addr_in[15]
  PIN addr_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END addr_in[16]
  PIN addr_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END addr_in[17]
  PIN addr_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END addr_in[18]
  PIN addr_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END addr_in[19]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 22.480 400.000 23.080 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 396.000 30.730 400.000 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 46.280 400.000 46.880 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 53.760 400.000 54.360 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 63.280 400.000 63.880 ;
    END
  END addr_in[9]
  PIN addr_to_core_mem[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END addr_to_core_mem[0]
  PIN addr_to_core_mem[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END addr_to_core_mem[10]
  PIN addr_to_core_mem[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 79.600 400.000 80.200 ;
    END
  END addr_to_core_mem[11]
  PIN addr_to_core_mem[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 396.000 77.650 400.000 ;
    END
  END addr_to_core_mem[12]
  PIN addr_to_core_mem[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 87.080 400.000 87.680 ;
    END
  END addr_to_core_mem[13]
  PIN addr_to_core_mem[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END addr_to_core_mem[14]
  PIN addr_to_core_mem[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END addr_to_core_mem[15]
  PIN addr_to_core_mem[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 396.000 97.890 400.000 ;
    END
  END addr_to_core_mem[16]
  PIN addr_to_core_mem[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END addr_to_core_mem[17]
  PIN addr_to_core_mem[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 396.000 106.170 400.000 ;
    END
  END addr_to_core_mem[18]
  PIN addr_to_core_mem[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 396.000 112.610 400.000 ;
    END
  END addr_to_core_mem[19]
  PIN addr_to_core_mem[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END addr_to_core_mem[1]
  PIN addr_to_core_mem[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 396.000 14.170 400.000 ;
    END
  END addr_to_core_mem[2]
  PIN addr_to_core_mem[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 396.000 22.450 400.000 ;
    END
  END addr_to_core_mem[3]
  PIN addr_to_core_mem[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END addr_to_core_mem[4]
  PIN addr_to_core_mem[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END addr_to_core_mem[5]
  PIN addr_to_core_mem[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 42.880 400.000 43.480 ;
    END
  END addr_to_core_mem[6]
  PIN addr_to_core_mem[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 48.320 400.000 48.920 ;
    END
  END addr_to_core_mem[7]
  PIN addr_to_core_mem[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 396.000 54.190 400.000 ;
    END
  END addr_to_core_mem[8]
  PIN addr_to_core_mem[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 64.640 400.000 65.240 ;
    END
  END addr_to_core_mem[9]
  PIN clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END clk
  PIN core0_data_print[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 396.000 2.210 400.000 ;
    END
  END core0_data_print[0]
  PIN core0_data_print[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END core0_data_print[10]
  PIN core0_data_print[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 396.000 64.310 400.000 ;
    END
  END core0_data_print[11]
  PIN core0_data_print[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END core0_data_print[12]
  PIN core0_data_print[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 396.000 82.710 400.000 ;
    END
  END core0_data_print[13]
  PIN core0_data_print[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 97.960 400.000 98.560 ;
    END
  END core0_data_print[14]
  PIN core0_data_print[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 108.840 400.000 109.440 ;
    END
  END core0_data_print[15]
  PIN core0_data_print[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 396.000 99.270 400.000 ;
    END
  END core0_data_print[16]
  PIN core0_data_print[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END core0_data_print[17]
  PIN core0_data_print[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END core0_data_print[18]
  PIN core0_data_print[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 396.000 114.450 400.000 ;
    END
  END core0_data_print[19]
  PIN core0_data_print[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 396.000 9.110 400.000 ;
    END
  END core0_data_print[1]
  PIN core0_data_print[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END core0_data_print[20]
  PIN core0_data_print[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 396.000 124.570 400.000 ;
    END
  END core0_data_print[21]
  PIN core0_data_print[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END core0_data_print[22]
  PIN core0_data_print[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END core0_data_print[23]
  PIN core0_data_print[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 157.120 400.000 157.720 ;
    END
  END core0_data_print[24]
  PIN core0_data_print[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END core0_data_print[25]
  PIN core0_data_print[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 165.960 400.000 166.560 ;
    END
  END core0_data_print[26]
  PIN core0_data_print[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END core0_data_print[27]
  PIN core0_data_print[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 396.000 164.590 400.000 ;
    END
  END core0_data_print[28]
  PIN core0_data_print[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END core0_data_print[29]
  PIN core0_data_print[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 12.960 400.000 13.560 ;
    END
  END core0_data_print[2]
  PIN core0_data_print[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 188.400 400.000 189.000 ;
    END
  END core0_data_print[30]
  PIN core0_data_print[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END core0_data_print[31]
  PIN core0_data_print[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 396.000 23.830 400.000 ;
    END
  END core0_data_print[3]
  PIN core0_data_print[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 24.520 400.000 25.120 ;
    END
  END core0_data_print[4]
  PIN core0_data_print[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END core0_data_print[5]
  PIN core0_data_print[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END core0_data_print[6]
  PIN core0_data_print[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END core0_data_print[7]
  PIN core0_data_print[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END core0_data_print[8]
  PIN core0_data_print[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END core0_data_print[9]
  PIN csb0_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 2.080 400.000 2.680 ;
    END
  END csb0_to_sram
  PIN data_out_to_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END data_out_to_core[0]
  PIN data_out_to_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 74.160 400.000 74.760 ;
    END
  END data_out_to_core[10]
  PIN data_out_to_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END data_out_to_core[11]
  PIN data_out_to_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 396.000 79.490 400.000 ;
    END
  END data_out_to_core[12]
  PIN data_out_to_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 89.120 400.000 89.720 ;
    END
  END data_out_to_core[13]
  PIN data_out_to_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 100.000 400.000 100.600 ;
    END
  END data_out_to_core[14]
  PIN data_out_to_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END data_out_to_core[15]
  PIN data_out_to_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 120.400 400.000 121.000 ;
    END
  END data_out_to_core[16]
  PIN data_out_to_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.240 400.000 129.840 ;
    END
  END data_out_to_core[17]
  PIN data_out_to_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END data_out_to_core[18]
  PIN data_out_to_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END data_out_to_core[19]
  PIN data_out_to_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 396.000 10.490 400.000 ;
    END
  END data_out_to_core[1]
  PIN data_out_to_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END data_out_to_core[20]
  PIN data_out_to_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END data_out_to_core[21]
  PIN data_out_to_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 396.000 136.070 400.000 ;
    END
  END data_out_to_core[22]
  PIN data_out_to_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 153.040 400.000 153.640 ;
    END
  END data_out_to_core[23]
  PIN data_out_to_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END data_out_to_core[24]
  PIN data_out_to_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END data_out_to_core[25]
  PIN data_out_to_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END data_out_to_core[26]
  PIN data_out_to_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 172.080 400.000 172.680 ;
    END
  END data_out_to_core[27]
  PIN data_out_to_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.920 400.000 181.520 ;
    END
  END data_out_to_core[28]
  PIN data_out_to_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 396.000 166.430 400.000 ;
    END
  END data_out_to_core[29]
  PIN data_out_to_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END data_out_to_core[2]
  PIN data_out_to_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 396.000 174.710 400.000 ;
    END
  END data_out_to_core[30]
  PIN data_out_to_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END data_out_to_core[31]
  PIN data_out_to_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END data_out_to_core[3]
  PIN data_out_to_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END data_out_to_core[4]
  PIN data_out_to_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 35.400 400.000 36.000 ;
    END
  END data_out_to_core[5]
  PIN data_out_to_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END data_out_to_core[6]
  PIN data_out_to_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 50.360 400.000 50.960 ;
    END
  END data_out_to_core[7]
  PIN data_out_to_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 55.800 400.000 56.400 ;
    END
  END data_out_to_core[8]
  PIN data_out_to_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END data_out_to_core[9]
  PIN data_to_core_mem[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END data_to_core_mem[0]
  PIN data_to_core_mem[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END data_to_core_mem[10]
  PIN data_to_core_mem[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END data_to_core_mem[11]
  PIN data_to_core_mem[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END data_to_core_mem[12]
  PIN data_to_core_mem[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END data_to_core_mem[13]
  PIN data_to_core_mem[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 102.040 400.000 102.640 ;
    END
  END data_to_core_mem[14]
  PIN data_to_core_mem[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 396.000 92.830 400.000 ;
    END
  END data_to_core_mem[15]
  PIN data_to_core_mem[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END data_to_core_mem[16]
  PIN data_to_core_mem[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 396.000 102.950 400.000 ;
    END
  END data_to_core_mem[17]
  PIN data_to_core_mem[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 396.000 107.550 400.000 ;
    END
  END data_to_core_mem[18]
  PIN data_to_core_mem[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END data_to_core_mem[19]
  PIN data_to_core_mem[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END data_to_core_mem[1]
  PIN data_to_core_mem[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END data_to_core_mem[20]
  PIN data_to_core_mem[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 396.000 126.410 400.000 ;
    END
  END data_to_core_mem[21]
  PIN data_to_core_mem[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END data_to_core_mem[22]
  PIN data_to_core_mem[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 396.000 142.970 400.000 ;
    END
  END data_to_core_mem[23]
  PIN data_to_core_mem[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 396.000 151.250 400.000 ;
    END
  END data_to_core_mem[24]
  PIN data_to_core_mem[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END data_to_core_mem[25]
  PIN data_to_core_mem[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END data_to_core_mem[26]
  PIN data_to_core_mem[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 396.000 159.530 400.000 ;
    END
  END data_to_core_mem[27]
  PIN data_to_core_mem[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END data_to_core_mem[28]
  PIN data_to_core_mem[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 184.320 400.000 184.920 ;
    END
  END data_to_core_mem[29]
  PIN data_to_core_mem[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 396.000 15.550 400.000 ;
    END
  END data_to_core_mem[2]
  PIN data_to_core_mem[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END data_to_core_mem[30]
  PIN data_to_core_mem[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END data_to_core_mem[31]
  PIN data_to_core_mem[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 17.040 400.000 17.640 ;
    END
  END data_to_core_mem[3]
  PIN data_to_core_mem[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END data_to_core_mem[4]
  PIN data_to_core_mem[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END data_to_core_mem[5]
  PIN data_to_core_mem[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END data_to_core_mem[6]
  PIN data_to_core_mem[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END data_to_core_mem[7]
  PIN data_to_core_mem[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END data_to_core_mem[8]
  PIN data_to_core_mem[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 66.680 400.000 67.280 ;
    END
  END data_to_core_mem[9]
  PIN din0_to_sram[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 396.000 4.050 400.000 ;
    END
  END din0_to_sram[0]
  PIN din0_to_sram[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END din0_to_sram[10]
  PIN din0_to_sram[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 396.000 65.690 400.000 ;
    END
  END din0_to_sram[11]
  PIN din0_to_sram[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END din0_to_sram[12]
  PIN din0_to_sram[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END din0_to_sram[13]
  PIN din0_to_sram[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 396.000 84.550 400.000 ;
    END
  END din0_to_sram[14]
  PIN din0_to_sram[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 110.880 400.000 111.480 ;
    END
  END din0_to_sram[15]
  PIN din0_to_sram[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 121.760 400.000 122.360 ;
    END
  END din0_to_sram[16]
  PIN din0_to_sram[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END din0_to_sram[17]
  PIN din0_to_sram[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 396.000 109.390 400.000 ;
    END
  END din0_to_sram[18]
  PIN din0_to_sram[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.160 400.000 142.760 ;
    END
  END din0_to_sram[19]
  PIN din0_to_sram[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 396.000 12.330 400.000 ;
    END
  END din0_to_sram[1]
  PIN din0_to_sram[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END din0_to_sram[20]
  PIN din0_to_sram[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END din0_to_sram[21]
  PIN din0_to_sram[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 396.000 137.910 400.000 ;
    END
  END din0_to_sram[22]
  PIN din0_to_sram[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END din0_to_sram[23]
  PIN din0_to_sram[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.160 400.000 159.760 ;
    END
  END din0_to_sram[24]
  PIN din0_to_sram[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 164.600 400.000 165.200 ;
    END
  END din0_to_sram[25]
  PIN din0_to_sram[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 396.000 158.150 400.000 ;
    END
  END din0_to_sram[26]
  PIN din0_to_sram[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 173.440 400.000 174.040 ;
    END
  END din0_to_sram[27]
  PIN din0_to_sram[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END din0_to_sram[28]
  PIN din0_to_sram[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 396.000 168.270 400.000 ;
    END
  END din0_to_sram[29]
  PIN din0_to_sram[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 396.000 17.390 400.000 ;
    END
  END din0_to_sram[2]
  PIN din0_to_sram[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END din0_to_sram[30]
  PIN din0_to_sram[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 396.000 177.930 400.000 ;
    END
  END din0_to_sram[31]
  PIN din0_to_sram[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END din0_to_sram[3]
  PIN din0_to_sram[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END din0_to_sram[4]
  PIN din0_to_sram[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END din0_to_sram[5]
  PIN din0_to_sram[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 396.000 39.010 400.000 ;
    END
  END din0_to_sram[6]
  PIN din0_to_sram[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END din0_to_sram[7]
  PIN din0_to_sram[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END din0_to_sram[8]
  PIN din0_to_sram[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.720 400.000 69.320 ;
    END
  END din0_to_sram[9]
  PIN dout0_to_sram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 396.000 5.430 400.000 ;
    END
  END dout0_to_sram[0]
  PIN dout0_to_sram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 396.000 61.090 400.000 ;
    END
  END dout0_to_sram[10]
  PIN dout0_to_sram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 396.000 67.530 400.000 ;
    END
  END dout0_to_sram[11]
  PIN dout0_to_sram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END dout0_to_sram[12]
  PIN dout0_to_sram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 90.480 400.000 91.080 ;
    END
  END dout0_to_sram[13]
  PIN dout0_to_sram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 396.000 85.930 400.000 ;
    END
  END dout0_to_sram[14]
  PIN dout0_to_sram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END dout0_to_sram[15]
  PIN dout0_to_sram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END dout0_to_sram[16]
  PIN dout0_to_sram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 131.280 400.000 131.880 ;
    END
  END dout0_to_sram[17]
  PIN dout0_to_sram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 134.680 400.000 135.280 ;
    END
  END dout0_to_sram[18]
  PIN dout0_to_sram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 396.000 116.290 400.000 ;
    END
  END dout0_to_sram[19]
  PIN dout0_to_sram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END dout0_to_sram[1]
  PIN dout0_to_sram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END dout0_to_sram[20]
  PIN dout0_to_sram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 396.000 127.790 400.000 ;
    END
  END dout0_to_sram[21]
  PIN dout0_to_sram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END dout0_to_sram[22]
  PIN dout0_to_sram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 155.080 400.000 155.680 ;
    END
  END dout0_to_sram[23]
  PIN dout0_to_sram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END dout0_to_sram[24]
  PIN dout0_to_sram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END dout0_to_sram[25]
  PIN dout0_to_sram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END dout0_to_sram[26]
  PIN dout0_to_sram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 175.480 400.000 176.080 ;
    END
  END dout0_to_sram[27]
  PIN dout0_to_sram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END dout0_to_sram[28]
  PIN dout0_to_sram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 186.360 400.000 186.960 ;
    END
  END dout0_to_sram[29]
  PIN dout0_to_sram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 396.000 19.230 400.000 ;
    END
  END dout0_to_sram[2]
  PIN dout0_to_sram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END dout0_to_sram[30]
  PIN dout0_to_sram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 396.000 179.770 400.000 ;
    END
  END dout0_to_sram[31]
  PIN dout0_to_sram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 396.000 25.670 400.000 ;
    END
  END dout0_to_sram[3]
  PIN dout0_to_sram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 25.880 400.000 26.480 ;
    END
  END dout0_to_sram[4]
  PIN dout0_to_sram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 37.440 400.000 38.040 ;
    END
  END dout0_to_sram[5]
  PIN dout0_to_sram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END dout0_to_sram[6]
  PIN dout0_to_sram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END dout0_to_sram[7]
  PIN dout0_to_sram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 57.840 400.000 58.440 ;
    END
  END dout0_to_sram[8]
  PIN dout0_to_sram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 396.000 59.250 400.000 ;
    END
  END dout0_to_sram[9]
  PIN is_loading_memory_into_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END is_loading_memory_into_core
  PIN is_ready_dataout_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END is_ready_dataout_core0
  PIN is_ready_print_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END is_ready_print_core0
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 396.000 350.430 400.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 350.240 400.000 350.840 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.520 4.000 348.120 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 365.200 400.000 365.800 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 367.240 400.000 367.840 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 396.000 365.610 400.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 396.000 367.450 400.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 378.120 400.000 378.720 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 396.000 69.370 400.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 81.640 400.000 82.240 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 92.520 400.000 93.120 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 396.000 87.770 400.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 396.000 94.210 400.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.800 400.000 124.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 136.720 400.000 137.320 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 396.000 119.510 400.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 396.000 129.630 400.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 396.000 139.750 400.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 396.000 144.810 400.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 160.520 400.000 161.120 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 396.000 161.370 400.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.240 400.000 197.840 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 199.280 400.000 199.880 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 396.000 194.950 400.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 203.360 400.000 203.960 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 396.000 205.070 400.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 396.000 206.450 400.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.240 400.000 214.840 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 396.000 214.730 400.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 225.120 400.000 225.720 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.160 400.000 227.760 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 396.000 27.510 400.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 396.000 223.470 400.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 236.000 400.000 236.600 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.920 400.000 249.520 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 38.800 400.000 39.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 396.000 241.870 400.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 256.400 400.000 257.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 261.840 400.000 262.440 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 263.880 400.000 264.480 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 396.000 268.550 400.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 396.000 271.770 400.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 273.400 400.000 274.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 396.000 278.670 400.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 396.000 292.010 400.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 396.000 293.850 400.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 396.000 297.070 400.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 396.000 300.290 400.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 289.720 400.000 290.320 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 396.000 45.910 400.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 291.760 400.000 292.360 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 298.560 400.000 299.160 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 396.000 315.470 400.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 323.040 400.000 323.640 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 396.000 320.530 400.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 396.000 56.030 400.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 396.000 326.970 400.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 335.960 400.000 336.560 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 339.360 400.000 339.960 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 396.000 345.370 400.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 346.840 400.000 347.440 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 352.280 400.000 352.880 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 396.000 355.490 400.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.720 400.000 358.320 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 359.760 400.000 360.360 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 76.200 400.000 76.800 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 374.720 400.000 375.320 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 376.080 400.000 376.680 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 396.000 375.730 400.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 381.520 400.000 382.120 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 396.000 385.850 400.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 396.000 390.910 400.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 396.000 394.130 400.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 396.480 400.000 397.080 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 396.000 89.150 400.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.920 400.000 113.520 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 138.760 400.000 139.360 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 396.000 131.010 400.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 396.000 156.310 400.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 168.000 400.000 168.600 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 177.520 400.000 178.120 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 191.800 400.000 192.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 201.320 400.000 201.920 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 396.000 198.170 400.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 396.000 201.390 400.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 19.080 400.000 19.680 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.720 400.000 205.320 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 208.800 400.000 209.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 396.000 208.290 400.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 219.680 400.000 220.280 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 396.000 211.510 400.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 27.920 400.000 28.520 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 396.000 224.850 400.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.040 400.000 238.640 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 243.480 400.000 244.080 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 396.000 231.750 400.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 247.560 400.000 248.160 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 396.000 236.810 400.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 396.000 32.570 400.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 250.960 400.000 251.560 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 253.000 400.000 253.600 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 396.000 246.930 400.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 396.000 253.370 400.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 396.000 256.590 400.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 396.000 261.650 400.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.920 400.000 266.520 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 396.000 270.390 400.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 269.320 400.000 269.920 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 44.920 400.000 45.520 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 274.760 400.000 275.360 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 396.000 280.050 400.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 396.000 285.110 400.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 282.240 400.000 282.840 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 286.320 400.000 286.920 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 396.000 303.510 400.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 396.000 47.290 400.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 396.000 307.190 400.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 302.640 400.000 303.240 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 304.680 400.000 305.280 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 308.080 400.000 308.680 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 396.000 316.850 400.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 396.000 325.590 400.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 396.000 328.810 400.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 396.000 333.870 400.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 396.000 337.090 400.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 341.400 400.000 342.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 343.440 400.000 344.040 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 396.000 347.210 400.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 6.160 400.000 6.760 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 354.320 400.000 354.920 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 368.600 400.000 369.200 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 396.000 370.670 400.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 396.000 373.890 400.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 396.000 377.570 400.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 396.000 378.950 400.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 383.560 400.000 384.160 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 396.000 382.170 400.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 396.000 384.010 400.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 396.000 70.750 400.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 387.640 400.000 388.240 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 396.000 389.070 400.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 391.040 400.000 391.640 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 396.000 395.970 400.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 396.000 399.190 400.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 94.560 400.000 95.160 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 396.000 90.990 400.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 114.960 400.000 115.560 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 125.840 400.000 126.440 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 396.000 111.230 400.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 144.200 400.000 144.800 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 396.000 132.850 400.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 396.000 141.130 400.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 396.000 146.190 400.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 396.000 153.090 400.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 178.880 400.000 179.480 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 182.960 400.000 183.560 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 396.000 20.610 400.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 190.440 400.000 191.040 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 195.880 400.000 196.480 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 396.000 191.270 400.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.280 400.000 216.880 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 396.000 216.570 400.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 396.000 219.790 400.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 229.200 400.000 229.800 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 29.960 400.000 30.560 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 396.000 226.690 400.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 396.000 228.530 400.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 396.000 233.130 400.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 396.000 234.970 400.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 396.000 33.950 400.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 396.000 243.250 400.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 254.360 400.000 254.960 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 396.000 248.310 400.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 396.000 258.430 400.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 396.000 265.330 400.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 267.280 400.000 267.880 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 396.000 273.610 400.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 396.000 40.850 400.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 276.800 400.000 277.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.840 400.000 279.440 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 396.000 286.950 400.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 396.000 49.130 400.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 293.120 400.000 293.720 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 396.000 310.410 400.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 396.000 312.250 400.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 310.120 400.000 310.720 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 313.520 400.000 314.120 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 318.960 400.000 319.560 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 396.000 318.690 400.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 396.000 321.910 400.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 396.000 57.410 400.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 330.520 400.000 331.120 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 396.000 330.650 400.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 396.000 338.930 400.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 344.800 400.000 345.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END la_oenb[9]
  PIN rd_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END rd_data_out[0]
  PIN rd_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 396.000 352.270 400.000 ;
    END
  END rd_data_out[100]
  PIN rd_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END rd_data_out[101]
  PIN rd_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 396.000 354.110 400.000 ;
    END
  END rd_data_out[102]
  PIN rd_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 355.680 400.000 356.280 ;
    END
  END rd_data_out[103]
  PIN rd_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 396.000 358.710 400.000 ;
    END
  END rd_data_out[104]
  PIN rd_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END rd_data_out[105]
  PIN rd_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 361.800 400.000 362.400 ;
    END
  END rd_data_out[106]
  PIN rd_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 396.000 362.390 400.000 ;
    END
  END rd_data_out[107]
  PIN rd_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END rd_data_out[108]
  PIN rd_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END rd_data_out[109]
  PIN rd_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END rd_data_out[10]
  PIN rd_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 396.000 363.770 400.000 ;
    END
  END rd_data_out[110]
  PIN rd_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END rd_data_out[111]
  PIN rd_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 372.680 400.000 373.280 ;
    END
  END rd_data_out[112]
  PIN rd_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END rd_data_out[113]
  PIN rd_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END rd_data_out[114]
  PIN rd_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END rd_data_out[115]
  PIN rd_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END rd_data_out[116]
  PIN rd_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 396.000 380.790 400.000 ;
    END
  END rd_data_out[117]
  PIN rd_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END rd_data_out[118]
  PIN rd_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 385.600 400.000 386.200 ;
    END
  END rd_data_out[119]
  PIN rd_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 396.000 72.590 400.000 ;
    END
  END rd_data_out[11]
  PIN rd_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END rd_data_out[120]
  PIN rd_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END rd_data_out[121]
  PIN rd_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 393.080 400.000 393.680 ;
    END
  END rd_data_out[122]
  PIN rd_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END rd_data_out[123]
  PIN rd_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 394.440 400.000 395.040 ;
    END
  END rd_data_out[124]
  PIN rd_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END rd_data_out[125]
  PIN rd_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END rd_data_out[126]
  PIN rd_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 398.520 400.000 399.120 ;
    END
  END rd_data_out[127]
  PIN rd_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 396.000 80.870 400.000 ;
    END
  END rd_data_out[12]
  PIN rd_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END rd_data_out[13]
  PIN rd_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END rd_data_out[14]
  PIN rd_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 116.320 400.000 116.920 ;
    END
  END rd_data_out[15]
  PIN rd_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END rd_data_out[16]
  PIN rd_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END rd_data_out[17]
  PIN rd_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END rd_data_out[18]
  PIN rd_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 146.240 400.000 146.840 ;
    END
  END rd_data_out[19]
  PIN rd_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END rd_data_out[1]
  PIN rd_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 396.000 121.350 400.000 ;
    END
  END rd_data_out[20]
  PIN rd_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 396.000 134.690 400.000 ;
    END
  END rd_data_out[21]
  PIN rd_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END rd_data_out[22]
  PIN rd_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END rd_data_out[23]
  PIN rd_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 396.000 154.470 400.000 ;
    END
  END rd_data_out[24]
  PIN rd_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END rd_data_out[25]
  PIN rd_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END rd_data_out[26]
  PIN rd_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END rd_data_out[27]
  PIN rd_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END rd_data_out[28]
  PIN rd_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END rd_data_out[29]
  PIN rd_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END rd_data_out[2]
  PIN rd_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END rd_data_out[30]
  PIN rd_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END rd_data_out[31]
  PIN rd_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END rd_data_out[32]
  PIN rd_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END rd_data_out[33]
  PIN rd_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END rd_data_out[34]
  PIN rd_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END rd_data_out[35]
  PIN rd_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END rd_data_out[36]
  PIN rd_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END rd_data_out[37]
  PIN rd_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 396.000 200.010 400.000 ;
    END
  END rd_data_out[38]
  PIN rd_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END rd_data_out[39]
  PIN rd_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END rd_data_out[3]
  PIN rd_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 396.000 203.230 400.000 ;
    END
  END rd_data_out[40]
  PIN rd_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END rd_data_out[41]
  PIN rd_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 206.760 400.000 207.360 ;
    END
  END rd_data_out[42]
  PIN rd_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.160 400.000 210.760 ;
    END
  END rd_data_out[43]
  PIN rd_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 217.640 400.000 218.240 ;
    END
  END rd_data_out[44]
  PIN rd_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.720 400.000 222.320 ;
    END
  END rd_data_out[45]
  PIN rd_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 396.000 213.350 400.000 ;
    END
  END rd_data_out[46]
  PIN rd_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 396.000 218.410 400.000 ;
    END
  END rd_data_out[47]
  PIN rd_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END rd_data_out[48]
  PIN rd_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 396.000 221.630 400.000 ;
    END
  END rd_data_out[49]
  PIN rd_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 32.000 400.000 32.600 ;
    END
  END rd_data_out[4]
  PIN rd_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END rd_data_out[50]
  PIN rd_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 232.600 400.000 233.200 ;
    END
  END rd_data_out[51]
  PIN rd_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END rd_data_out[52]
  PIN rd_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END rd_data_out[53]
  PIN rd_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 241.440 400.000 242.040 ;
    END
  END rd_data_out[54]
  PIN rd_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END rd_data_out[55]
  PIN rd_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END rd_data_out[56]
  PIN rd_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END rd_data_out[57]
  PIN rd_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END rd_data_out[58]
  PIN rd_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 396.000 238.190 400.000 ;
    END
  END rd_data_out[59]
  PIN rd_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 396.000 35.790 400.000 ;
    END
  END rd_data_out[5]
  PIN rd_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END rd_data_out[60]
  PIN rd_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END rd_data_out[61]
  PIN rd_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 396.000 250.150 400.000 ;
    END
  END rd_data_out[62]
  PIN rd_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 396.000 251.990 400.000 ;
    END
  END rd_data_out[63]
  PIN rd_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 396.000 255.210 400.000 ;
    END
  END rd_data_out[64]
  PIN rd_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END rd_data_out[65]
  PIN rd_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END rd_data_out[66]
  PIN rd_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END rd_data_out[67]
  PIN rd_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END rd_data_out[68]
  PIN rd_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 271.360 400.000 271.960 ;
    END
  END rd_data_out[69]
  PIN rd_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END rd_data_out[6]
  PIN rd_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 396.000 274.990 400.000 ;
    END
  END rd_data_out[70]
  PIN rd_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END rd_data_out[71]
  PIN rd_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END rd_data_out[72]
  PIN rd_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END rd_data_out[73]
  PIN rd_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 396.000 288.790 400.000 ;
    END
  END rd_data_out[74]
  PIN rd_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END rd_data_out[75]
  PIN rd_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 396.000 295.230 400.000 ;
    END
  END rd_data_out[76]
  PIN rd_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 284.280 400.000 284.880 ;
    END
  END rd_data_out[77]
  PIN rd_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 396.000 302.130 400.000 ;
    END
  END rd_data_out[78]
  PIN rd_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END rd_data_out[79]
  PIN rd_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 51.720 400.000 52.320 ;
    END
  END rd_data_out[7]
  PIN rd_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END rd_data_out[80]
  PIN rd_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 295.160 400.000 295.760 ;
    END
  END rd_data_out[81]
  PIN rd_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END rd_data_out[82]
  PIN rd_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 396.000 313.630 400.000 ;
    END
  END rd_data_out[83]
  PIN rd_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END rd_data_out[84]
  PIN rd_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 311.480 400.000 312.080 ;
    END
  END rd_data_out[85]
  PIN rd_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 315.560 400.000 316.160 ;
    END
  END rd_data_out[86]
  PIN rd_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END rd_data_out[87]
  PIN rd_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END rd_data_out[88]
  PIN rd_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 326.440 400.000 327.040 ;
    END
  END rd_data_out[89]
  PIN rd_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END rd_data_out[8]
  PIN rd_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END rd_data_out[90]
  PIN rd_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 331.880 400.000 332.480 ;
    END
  END rd_data_out[91]
  PIN rd_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END rd_data_out[92]
  PIN rd_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.920 400.000 334.520 ;
    END
  END rd_data_out[93]
  PIN rd_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 396.000 335.710 400.000 ;
    END
  END rd_data_out[94]
  PIN rd_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END rd_data_out[95]
  PIN rd_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 396.000 340.310 400.000 ;
    END
  END rd_data_out[96]
  PIN rd_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 396.000 343.990 400.000 ;
    END
  END rd_data_out[97]
  PIN rd_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END rd_data_out[98]
  PIN rd_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END rd_data_out[99]
  PIN rd_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END rd_data_out[9]
  PIN read_enable_to_Elpis
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END read_enable_to_Elpis
  PIN read_interactive_req_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END read_interactive_req_core0
  PIN read_value_to_Elpis[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 396.000 7.270 400.000 ;
    END
  END read_value_to_Elpis[0]
  PIN read_value_to_Elpis[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END read_value_to_Elpis[10]
  PIN read_value_to_Elpis[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END read_value_to_Elpis[11]
  PIN read_value_to_Elpis[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END read_value_to_Elpis[12]
  PIN read_value_to_Elpis[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END read_value_to_Elpis[13]
  PIN read_value_to_Elpis[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 103.400 400.000 104.000 ;
    END
  END read_value_to_Elpis[14]
  PIN read_value_to_Elpis[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END read_value_to_Elpis[15]
  PIN read_value_to_Elpis[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 396.000 101.110 400.000 ;
    END
  END read_value_to_Elpis[16]
  PIN read_value_to_Elpis[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END read_value_to_Elpis[17]
  PIN read_value_to_Elpis[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END read_value_to_Elpis[18]
  PIN read_value_to_Elpis[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 147.600 400.000 148.200 ;
    END
  END read_value_to_Elpis[19]
  PIN read_value_to_Elpis[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END read_value_to_Elpis[1]
  PIN read_value_to_Elpis[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END read_value_to_Elpis[20]
  PIN read_value_to_Elpis[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 149.640 400.000 150.240 ;
    END
  END read_value_to_Elpis[21]
  PIN read_value_to_Elpis[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END read_value_to_Elpis[22]
  PIN read_value_to_Elpis[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 396.000 148.030 400.000 ;
    END
  END read_value_to_Elpis[23]
  PIN read_value_to_Elpis[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END read_value_to_Elpis[24]
  PIN read_value_to_Elpis[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END read_value_to_Elpis[25]
  PIN read_value_to_Elpis[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END read_value_to_Elpis[26]
  PIN read_value_to_Elpis[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END read_value_to_Elpis[27]
  PIN read_value_to_Elpis[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END read_value_to_Elpis[28]
  PIN read_value_to_Elpis[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 396.000 169.650 400.000 ;
    END
  END read_value_to_Elpis[29]
  PIN read_value_to_Elpis[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END read_value_to_Elpis[2]
  PIN read_value_to_Elpis[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END read_value_to_Elpis[30]
  PIN read_value_to_Elpis[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 396.000 181.610 400.000 ;
    END
  END read_value_to_Elpis[31]
  PIN read_value_to_Elpis[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END read_value_to_Elpis[3]
  PIN read_value_to_Elpis[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 33.360 400.000 33.960 ;
    END
  END read_value_to_Elpis[4]
  PIN read_value_to_Elpis[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 40.840 400.000 41.440 ;
    END
  END read_value_to_Elpis[5]
  PIN read_value_to_Elpis[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 396.000 42.690 400.000 ;
    END
  END read_value_to_Elpis[6]
  PIN read_value_to_Elpis[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END read_value_to_Elpis[7]
  PIN read_value_to_Elpis[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END read_value_to_Elpis[8]
  PIN read_value_to_Elpis[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 70.080 400.000 70.680 ;
    END
  END read_value_to_Elpis[9]
  PIN ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END ready
  PIN req_out_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END req_out_core0
  PIN requested
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END requested
  PIN reset_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END reset_core
  PIN reset_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END reset_mem_req
  PIN rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END rst
  PIN spare_wen0_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 4.120 400.000 4.720 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_rst_i
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 7.520 400.000 8.120 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 396.000 74.430 400.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 83.000 400.000 83.600 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 396.000 96.050 400.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 396.000 104.330 400.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 396.000 149.410 400.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.040 400.000 170.640 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 396.000 171.490 400.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 15.000 400.000 15.600 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 396.000 176.550 400.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 396.000 182.990 400.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 396.000 37.630 400.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 396.000 50.970 400.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 59.200 400.000 59.800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END wbs_dat_o[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END we
  PIN we_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 0.720 400.000 1.320 ;
    END
  END we_to_sram
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END wr_data[0]
  PIN wr_data[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 348.880 400.000 349.480 ;
    END
  END wr_data[100]
  PIN wr_data[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END wr_data[101]
  PIN wr_data[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END wr_data[102]
  PIN wr_data[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 396.000 357.330 400.000 ;
    END
  END wr_data[103]
  PIN wr_data[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END wr_data[104]
  PIN wr_data[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 396.000 360.550 400.000 ;
    END
  END wr_data[105]
  PIN wr_data[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 363.160 400.000 363.760 ;
    END
  END wr_data[106]
  PIN wr_data[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END wr_data[107]
  PIN wr_data[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END wr_data[108]
  PIN wr_data[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END wr_data[109]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wr_data[10]
  PIN wr_data[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 370.640 400.000 371.240 ;
    END
  END wr_data[110]
  PIN wr_data[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END wr_data[111]
  PIN wr_data[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 396.000 368.830 400.000 ;
    END
  END wr_data[112]
  PIN wr_data[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 396.000 372.510 400.000 ;
    END
  END wr_data[113]
  PIN wr_data[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END wr_data[114]
  PIN wr_data[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END wr_data[115]
  PIN wr_data[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 380.160 400.000 380.760 ;
    END
  END wr_data[116]
  PIN wr_data[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END wr_data[117]
  PIN wr_data[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END wr_data[118]
  PIN wr_data[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END wr_data[119]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wr_data[11]
  PIN wr_data[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 396.000 387.230 400.000 ;
    END
  END wr_data[120]
  PIN wr_data[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 389.000 400.000 389.600 ;
    END
  END wr_data[121]
  PIN wr_data[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 396.000 392.290 400.000 ;
    END
  END wr_data[122]
  PIN wr_data[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END wr_data[123]
  PIN wr_data[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 396.000 397.350 400.000 ;
    END
  END wr_data[124]
  PIN wr_data[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END wr_data[125]
  PIN wr_data[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END wr_data[126]
  PIN wr_data[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END wr_data[127]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END wr_data[12]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END wr_data[13]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END wr_data[14]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 118.360 400.000 118.960 ;
    END
  END wr_data[15]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wr_data[16]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wr_data[17]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 140.120 400.000 140.720 ;
    END
  END wr_data[18]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 396.000 117.670 400.000 ;
    END
  END wr_data[19]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 11.600 400.000 12.200 ;
    END
  END wr_data[1]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 396.000 122.730 400.000 ;
    END
  END wr_data[20]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 151.680 400.000 152.280 ;
    END
  END wr_data[21]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END wr_data[22]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END wr_data[23]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 162.560 400.000 163.160 ;
    END
  END wr_data[24]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END wr_data[25]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END wr_data[26]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 396.000 163.210 400.000 ;
    END
  END wr_data[27]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END wr_data[28]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 396.000 172.870 400.000 ;
    END
  END wr_data[29]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wr_data[2]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wr_data[30]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 396.000 184.830 400.000 ;
    END
  END wr_data[31]
  PIN wr_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 396.000 186.670 400.000 ;
    END
  END wr_data[32]
  PIN wr_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.840 400.000 194.440 ;
    END
  END wr_data[33]
  PIN wr_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 396.000 188.050 400.000 ;
    END
  END wr_data[34]
  PIN wr_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 396.000 189.890 400.000 ;
    END
  END wr_data[35]
  PIN wr_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 396.000 193.110 400.000 ;
    END
  END wr_data[36]
  PIN wr_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 396.000 196.330 400.000 ;
    END
  END wr_data[37]
  PIN wr_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END wr_data[38]
  PIN wr_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END wr_data[39]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END wr_data[3]
  PIN wr_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END wr_data[40]
  PIN wr_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wr_data[41]
  PIN wr_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END wr_data[42]
  PIN wr_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 212.200 400.000 212.800 ;
    END
  END wr_data[43]
  PIN wr_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END wr_data[44]
  PIN wr_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 396.000 210.130 400.000 ;
    END
  END wr_data[45]
  PIN wr_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 223.080 400.000 223.680 ;
    END
  END wr_data[46]
  PIN wr_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END wr_data[47]
  PIN wr_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END wr_data[48]
  PIN wr_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END wr_data[49]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END wr_data[4]
  PIN wr_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 230.560 400.000 231.160 ;
    END
  END wr_data[50]
  PIN wr_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 234.640 400.000 235.240 ;
    END
  END wr_data[51]
  PIN wr_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 396.000 229.910 400.000 ;
    END
  END wr_data[52]
  PIN wr_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 240.080 400.000 240.680 ;
    END
  END wr_data[53]
  PIN wr_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END wr_data[54]
  PIN wr_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wr_data[55]
  PIN wr_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 245.520 400.000 246.120 ;
    END
  END wr_data[56]
  PIN wr_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END wr_data[57]
  PIN wr_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END wr_data[58]
  PIN wr_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 396.000 240.030 400.000 ;
    END
  END wr_data[59]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END wr_data[5]
  PIN wr_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 396.000 245.090 400.000 ;
    END
  END wr_data[60]
  PIN wr_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END wr_data[61]
  PIN wr_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 258.440 400.000 259.040 ;
    END
  END wr_data[62]
  PIN wr_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END wr_data[63]
  PIN wr_data[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 260.480 400.000 261.080 ;
    END
  END wr_data[64]
  PIN wr_data[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 396.000 260.270 400.000 ;
    END
  END wr_data[65]
  PIN wr_data[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 396.000 263.490 400.000 ;
    END
  END wr_data[66]
  PIN wr_data[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 396.000 266.710 400.000 ;
    END
  END wr_data[67]
  PIN wr_data[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END wr_data[68]
  PIN wr_data[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END wr_data[69]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wr_data[6]
  PIN wr_data[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 396.000 276.830 400.000 ;
    END
  END wr_data[70]
  PIN wr_data[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 396.000 281.890 400.000 ;
    END
  END wr_data[71]
  PIN wr_data[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 396.000 283.730 400.000 ;
    END
  END wr_data[72]
  PIN wr_data[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wr_data[73]
  PIN wr_data[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 396.000 290.170 400.000 ;
    END
  END wr_data[74]
  PIN wr_data[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 280.200 400.000 280.800 ;
    END
  END wr_data[75]
  PIN wr_data[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END wr_data[76]
  PIN wr_data[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 396.000 298.450 400.000 ;
    END
  END wr_data[77]
  PIN wr_data[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 287.680 400.000 288.280 ;
    END
  END wr_data[78]
  PIN wr_data[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 396.000 305.350 400.000 ;
    END
  END wr_data[79]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 396.000 52.350 400.000 ;
    END
  END wr_data[7]
  PIN wr_data[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 396.000 308.570 400.000 ;
    END
  END wr_data[80]
  PIN wr_data[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 297.200 400.000 297.800 ;
    END
  END wr_data[81]
  PIN wr_data[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 300.600 400.000 301.200 ;
    END
  END wr_data[82]
  PIN wr_data[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wr_data[83]
  PIN wr_data[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.040 400.000 306.640 ;
    END
  END wr_data[84]
  PIN wr_data[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END wr_data[85]
  PIN wr_data[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 317.600 400.000 318.200 ;
    END
  END wr_data[86]
  PIN wr_data[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.000 400.000 321.600 ;
    END
  END wr_data[87]
  PIN wr_data[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 324.400 400.000 325.000 ;
    END
  END wr_data[88]
  PIN wr_data[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END wr_data[89]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wr_data[8]
  PIN wr_data[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 328.480 400.000 329.080 ;
    END
  END wr_data[90]
  PIN wr_data[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 396.000 323.750 400.000 ;
    END
  END wr_data[91]
  PIN wr_data[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END wr_data[92]
  PIN wr_data[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 396.000 332.030 400.000 ;
    END
  END wr_data[93]
  PIN wr_data[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wr_data[94]
  PIN wr_data[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 337.320 400.000 337.920 ;
    END
  END wr_data[95]
  PIN wr_data[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 396.000 342.150 400.000 ;
    END
  END wr_data[96]
  PIN wr_data[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wr_data[97]
  PIN wr_data[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END wr_data[98]
  PIN wr_data[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 396.000 349.050 400.000 ;
    END
  END wr_data[99]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wr_data[9]
  OBS
      LAYER li1 ;
        RECT 4.745 9.945 396.835 394.655 ;
      LAYER met1 ;
        RECT 0.530 1.060 399.210 394.700 ;
      LAYER met2 ;
        RECT 1.110 395.720 1.650 399.005 ;
        RECT 2.490 395.720 3.490 399.005 ;
        RECT 4.330 395.720 4.870 399.005 ;
        RECT 5.710 395.720 6.710 399.005 ;
        RECT 7.550 395.720 8.550 399.005 ;
        RECT 9.390 395.720 9.930 399.005 ;
        RECT 10.770 395.720 11.770 399.005 ;
        RECT 12.610 395.720 13.610 399.005 ;
        RECT 14.450 395.720 14.990 399.005 ;
        RECT 15.830 395.720 16.830 399.005 ;
        RECT 17.670 395.720 18.670 399.005 ;
        RECT 19.510 395.720 20.050 399.005 ;
        RECT 20.890 395.720 21.890 399.005 ;
        RECT 22.730 395.720 23.270 399.005 ;
        RECT 24.110 395.720 25.110 399.005 ;
        RECT 25.950 395.720 26.950 399.005 ;
        RECT 27.790 395.720 28.330 399.005 ;
        RECT 29.170 395.720 30.170 399.005 ;
        RECT 31.010 395.720 32.010 399.005 ;
        RECT 32.850 395.720 33.390 399.005 ;
        RECT 34.230 395.720 35.230 399.005 ;
        RECT 36.070 395.720 37.070 399.005 ;
        RECT 37.910 395.720 38.450 399.005 ;
        RECT 39.290 395.720 40.290 399.005 ;
        RECT 41.130 395.720 42.130 399.005 ;
        RECT 42.970 395.720 43.510 399.005 ;
        RECT 44.350 395.720 45.350 399.005 ;
        RECT 46.190 395.720 46.730 399.005 ;
        RECT 47.570 395.720 48.570 399.005 ;
        RECT 49.410 395.720 50.410 399.005 ;
        RECT 51.250 395.720 51.790 399.005 ;
        RECT 52.630 395.720 53.630 399.005 ;
        RECT 54.470 395.720 55.470 399.005 ;
        RECT 56.310 395.720 56.850 399.005 ;
        RECT 57.690 395.720 58.690 399.005 ;
        RECT 59.530 395.720 60.530 399.005 ;
        RECT 61.370 395.720 61.910 399.005 ;
        RECT 62.750 395.720 63.750 399.005 ;
        RECT 64.590 395.720 65.130 399.005 ;
        RECT 65.970 395.720 66.970 399.005 ;
        RECT 67.810 395.720 68.810 399.005 ;
        RECT 69.650 395.720 70.190 399.005 ;
        RECT 71.030 395.720 72.030 399.005 ;
        RECT 72.870 395.720 73.870 399.005 ;
        RECT 74.710 395.720 75.250 399.005 ;
        RECT 76.090 395.720 77.090 399.005 ;
        RECT 77.930 395.720 78.930 399.005 ;
        RECT 79.770 395.720 80.310 399.005 ;
        RECT 81.150 395.720 82.150 399.005 ;
        RECT 82.990 395.720 83.990 399.005 ;
        RECT 84.830 395.720 85.370 399.005 ;
        RECT 86.210 395.720 87.210 399.005 ;
        RECT 88.050 395.720 88.590 399.005 ;
        RECT 89.430 395.720 90.430 399.005 ;
        RECT 91.270 395.720 92.270 399.005 ;
        RECT 93.110 395.720 93.650 399.005 ;
        RECT 94.490 395.720 95.490 399.005 ;
        RECT 96.330 395.720 97.330 399.005 ;
        RECT 98.170 395.720 98.710 399.005 ;
        RECT 99.550 395.720 100.550 399.005 ;
        RECT 101.390 395.720 102.390 399.005 ;
        RECT 103.230 395.720 103.770 399.005 ;
        RECT 104.610 395.720 105.610 399.005 ;
        RECT 106.450 395.720 106.990 399.005 ;
        RECT 107.830 395.720 108.830 399.005 ;
        RECT 109.670 395.720 110.670 399.005 ;
        RECT 111.510 395.720 112.050 399.005 ;
        RECT 112.890 395.720 113.890 399.005 ;
        RECT 114.730 395.720 115.730 399.005 ;
        RECT 116.570 395.720 117.110 399.005 ;
        RECT 117.950 395.720 118.950 399.005 ;
        RECT 119.790 395.720 120.790 399.005 ;
        RECT 121.630 395.720 122.170 399.005 ;
        RECT 123.010 395.720 124.010 399.005 ;
        RECT 124.850 395.720 125.850 399.005 ;
        RECT 126.690 395.720 127.230 399.005 ;
        RECT 128.070 395.720 129.070 399.005 ;
        RECT 129.910 395.720 130.450 399.005 ;
        RECT 131.290 395.720 132.290 399.005 ;
        RECT 133.130 395.720 134.130 399.005 ;
        RECT 134.970 395.720 135.510 399.005 ;
        RECT 136.350 395.720 137.350 399.005 ;
        RECT 138.190 395.720 139.190 399.005 ;
        RECT 140.030 395.720 140.570 399.005 ;
        RECT 141.410 395.720 142.410 399.005 ;
        RECT 143.250 395.720 144.250 399.005 ;
        RECT 145.090 395.720 145.630 399.005 ;
        RECT 146.470 395.720 147.470 399.005 ;
        RECT 148.310 395.720 148.850 399.005 ;
        RECT 149.690 395.720 150.690 399.005 ;
        RECT 151.530 395.720 152.530 399.005 ;
        RECT 153.370 395.720 153.910 399.005 ;
        RECT 154.750 395.720 155.750 399.005 ;
        RECT 156.590 395.720 157.590 399.005 ;
        RECT 158.430 395.720 158.970 399.005 ;
        RECT 159.810 395.720 160.810 399.005 ;
        RECT 161.650 395.720 162.650 399.005 ;
        RECT 163.490 395.720 164.030 399.005 ;
        RECT 164.870 395.720 165.870 399.005 ;
        RECT 166.710 395.720 167.710 399.005 ;
        RECT 168.550 395.720 169.090 399.005 ;
        RECT 169.930 395.720 170.930 399.005 ;
        RECT 171.770 395.720 172.310 399.005 ;
        RECT 173.150 395.720 174.150 399.005 ;
        RECT 174.990 395.720 175.990 399.005 ;
        RECT 176.830 395.720 177.370 399.005 ;
        RECT 178.210 395.720 179.210 399.005 ;
        RECT 180.050 395.720 181.050 399.005 ;
        RECT 181.890 395.720 182.430 399.005 ;
        RECT 183.270 395.720 184.270 399.005 ;
        RECT 185.110 395.720 186.110 399.005 ;
        RECT 186.950 395.720 187.490 399.005 ;
        RECT 188.330 395.720 189.330 399.005 ;
        RECT 190.170 395.720 190.710 399.005 ;
        RECT 191.550 395.720 192.550 399.005 ;
        RECT 193.390 395.720 194.390 399.005 ;
        RECT 195.230 395.720 195.770 399.005 ;
        RECT 196.610 395.720 197.610 399.005 ;
        RECT 198.450 395.720 199.450 399.005 ;
        RECT 200.290 395.720 200.830 399.005 ;
        RECT 201.670 395.720 202.670 399.005 ;
        RECT 203.510 395.720 204.510 399.005 ;
        RECT 205.350 395.720 205.890 399.005 ;
        RECT 206.730 395.720 207.730 399.005 ;
        RECT 208.570 395.720 209.570 399.005 ;
        RECT 210.410 395.720 210.950 399.005 ;
        RECT 211.790 395.720 212.790 399.005 ;
        RECT 213.630 395.720 214.170 399.005 ;
        RECT 215.010 395.720 216.010 399.005 ;
        RECT 216.850 395.720 217.850 399.005 ;
        RECT 218.690 395.720 219.230 399.005 ;
        RECT 220.070 395.720 221.070 399.005 ;
        RECT 221.910 395.720 222.910 399.005 ;
        RECT 223.750 395.720 224.290 399.005 ;
        RECT 225.130 395.720 226.130 399.005 ;
        RECT 226.970 395.720 227.970 399.005 ;
        RECT 228.810 395.720 229.350 399.005 ;
        RECT 230.190 395.720 231.190 399.005 ;
        RECT 232.030 395.720 232.570 399.005 ;
        RECT 233.410 395.720 234.410 399.005 ;
        RECT 235.250 395.720 236.250 399.005 ;
        RECT 237.090 395.720 237.630 399.005 ;
        RECT 238.470 395.720 239.470 399.005 ;
        RECT 240.310 395.720 241.310 399.005 ;
        RECT 242.150 395.720 242.690 399.005 ;
        RECT 243.530 395.720 244.530 399.005 ;
        RECT 245.370 395.720 246.370 399.005 ;
        RECT 247.210 395.720 247.750 399.005 ;
        RECT 248.590 395.720 249.590 399.005 ;
        RECT 250.430 395.720 251.430 399.005 ;
        RECT 252.270 395.720 252.810 399.005 ;
        RECT 253.650 395.720 254.650 399.005 ;
        RECT 255.490 395.720 256.030 399.005 ;
        RECT 256.870 395.720 257.870 399.005 ;
        RECT 258.710 395.720 259.710 399.005 ;
        RECT 260.550 395.720 261.090 399.005 ;
        RECT 261.930 395.720 262.930 399.005 ;
        RECT 263.770 395.720 264.770 399.005 ;
        RECT 265.610 395.720 266.150 399.005 ;
        RECT 266.990 395.720 267.990 399.005 ;
        RECT 268.830 395.720 269.830 399.005 ;
        RECT 270.670 395.720 271.210 399.005 ;
        RECT 272.050 395.720 273.050 399.005 ;
        RECT 273.890 395.720 274.430 399.005 ;
        RECT 275.270 395.720 276.270 399.005 ;
        RECT 277.110 395.720 278.110 399.005 ;
        RECT 278.950 395.720 279.490 399.005 ;
        RECT 280.330 395.720 281.330 399.005 ;
        RECT 282.170 395.720 283.170 399.005 ;
        RECT 284.010 395.720 284.550 399.005 ;
        RECT 285.390 395.720 286.390 399.005 ;
        RECT 287.230 395.720 288.230 399.005 ;
        RECT 289.070 395.720 289.610 399.005 ;
        RECT 290.450 395.720 291.450 399.005 ;
        RECT 292.290 395.720 293.290 399.005 ;
        RECT 294.130 395.720 294.670 399.005 ;
        RECT 295.510 395.720 296.510 399.005 ;
        RECT 297.350 395.720 297.890 399.005 ;
        RECT 298.730 395.720 299.730 399.005 ;
        RECT 300.570 395.720 301.570 399.005 ;
        RECT 302.410 395.720 302.950 399.005 ;
        RECT 303.790 395.720 304.790 399.005 ;
        RECT 305.630 395.720 306.630 399.005 ;
        RECT 307.470 395.720 308.010 399.005 ;
        RECT 308.850 395.720 309.850 399.005 ;
        RECT 310.690 395.720 311.690 399.005 ;
        RECT 312.530 395.720 313.070 399.005 ;
        RECT 313.910 395.720 314.910 399.005 ;
        RECT 315.750 395.720 316.290 399.005 ;
        RECT 317.130 395.720 318.130 399.005 ;
        RECT 318.970 395.720 319.970 399.005 ;
        RECT 320.810 395.720 321.350 399.005 ;
        RECT 322.190 395.720 323.190 399.005 ;
        RECT 324.030 395.720 325.030 399.005 ;
        RECT 325.870 395.720 326.410 399.005 ;
        RECT 327.250 395.720 328.250 399.005 ;
        RECT 329.090 395.720 330.090 399.005 ;
        RECT 330.930 395.720 331.470 399.005 ;
        RECT 332.310 395.720 333.310 399.005 ;
        RECT 334.150 395.720 335.150 399.005 ;
        RECT 335.990 395.720 336.530 399.005 ;
        RECT 337.370 395.720 338.370 399.005 ;
        RECT 339.210 395.720 339.750 399.005 ;
        RECT 340.590 395.720 341.590 399.005 ;
        RECT 342.430 395.720 343.430 399.005 ;
        RECT 344.270 395.720 344.810 399.005 ;
        RECT 345.650 395.720 346.650 399.005 ;
        RECT 347.490 395.720 348.490 399.005 ;
        RECT 349.330 395.720 349.870 399.005 ;
        RECT 350.710 395.720 351.710 399.005 ;
        RECT 352.550 395.720 353.550 399.005 ;
        RECT 354.390 395.720 354.930 399.005 ;
        RECT 355.770 395.720 356.770 399.005 ;
        RECT 357.610 395.720 358.150 399.005 ;
        RECT 358.990 395.720 359.990 399.005 ;
        RECT 360.830 395.720 361.830 399.005 ;
        RECT 362.670 395.720 363.210 399.005 ;
        RECT 364.050 395.720 365.050 399.005 ;
        RECT 365.890 395.720 366.890 399.005 ;
        RECT 367.730 395.720 368.270 399.005 ;
        RECT 369.110 395.720 370.110 399.005 ;
        RECT 370.950 395.720 371.950 399.005 ;
        RECT 372.790 395.720 373.330 399.005 ;
        RECT 374.170 395.720 375.170 399.005 ;
        RECT 376.010 395.720 377.010 399.005 ;
        RECT 377.850 395.720 378.390 399.005 ;
        RECT 379.230 395.720 380.230 399.005 ;
        RECT 381.070 395.720 381.610 399.005 ;
        RECT 382.450 395.720 383.450 399.005 ;
        RECT 384.290 395.720 385.290 399.005 ;
        RECT 386.130 395.720 386.670 399.005 ;
        RECT 387.510 395.720 388.510 399.005 ;
        RECT 389.350 395.720 390.350 399.005 ;
        RECT 391.190 395.720 391.730 399.005 ;
        RECT 392.570 395.720 393.570 399.005 ;
        RECT 394.410 395.720 395.410 399.005 ;
        RECT 396.250 395.720 396.790 399.005 ;
        RECT 397.630 395.720 398.630 399.005 ;
        RECT 0.560 4.280 399.180 395.720 ;
        RECT 1.110 0.835 1.650 4.280 ;
        RECT 2.490 0.835 3.030 4.280 ;
        RECT 3.870 0.835 4.870 4.280 ;
        RECT 5.710 0.835 6.250 4.280 ;
        RECT 7.090 0.835 8.090 4.280 ;
        RECT 8.930 0.835 9.470 4.280 ;
        RECT 10.310 0.835 11.310 4.280 ;
        RECT 12.150 0.835 12.690 4.280 ;
        RECT 13.530 0.835 14.530 4.280 ;
        RECT 15.370 0.835 15.910 4.280 ;
        RECT 16.750 0.835 17.750 4.280 ;
        RECT 18.590 0.835 19.130 4.280 ;
        RECT 19.970 0.835 20.970 4.280 ;
        RECT 21.810 0.835 22.350 4.280 ;
        RECT 23.190 0.835 24.190 4.280 ;
        RECT 25.030 0.835 25.570 4.280 ;
        RECT 26.410 0.835 27.410 4.280 ;
        RECT 28.250 0.835 28.790 4.280 ;
        RECT 29.630 0.835 30.630 4.280 ;
        RECT 31.470 0.835 32.010 4.280 ;
        RECT 32.850 0.835 33.850 4.280 ;
        RECT 34.690 0.835 35.230 4.280 ;
        RECT 36.070 0.835 37.070 4.280 ;
        RECT 37.910 0.835 38.450 4.280 ;
        RECT 39.290 0.835 40.290 4.280 ;
        RECT 41.130 0.835 41.670 4.280 ;
        RECT 42.510 0.835 43.050 4.280 ;
        RECT 43.890 0.835 44.890 4.280 ;
        RECT 45.730 0.835 46.270 4.280 ;
        RECT 47.110 0.835 48.110 4.280 ;
        RECT 48.950 0.835 49.490 4.280 ;
        RECT 50.330 0.835 51.330 4.280 ;
        RECT 52.170 0.835 52.710 4.280 ;
        RECT 53.550 0.835 54.550 4.280 ;
        RECT 55.390 0.835 55.930 4.280 ;
        RECT 56.770 0.835 57.770 4.280 ;
        RECT 58.610 0.835 59.150 4.280 ;
        RECT 59.990 0.835 60.990 4.280 ;
        RECT 61.830 0.835 62.370 4.280 ;
        RECT 63.210 0.835 64.210 4.280 ;
        RECT 65.050 0.835 65.590 4.280 ;
        RECT 66.430 0.835 67.430 4.280 ;
        RECT 68.270 0.835 68.810 4.280 ;
        RECT 69.650 0.835 70.650 4.280 ;
        RECT 71.490 0.835 72.030 4.280 ;
        RECT 72.870 0.835 73.870 4.280 ;
        RECT 74.710 0.835 75.250 4.280 ;
        RECT 76.090 0.835 77.090 4.280 ;
        RECT 77.930 0.835 78.470 4.280 ;
        RECT 79.310 0.835 80.310 4.280 ;
        RECT 81.150 0.835 81.690 4.280 ;
        RECT 82.530 0.835 83.070 4.280 ;
        RECT 83.910 0.835 84.910 4.280 ;
        RECT 85.750 0.835 86.290 4.280 ;
        RECT 87.130 0.835 88.130 4.280 ;
        RECT 88.970 0.835 89.510 4.280 ;
        RECT 90.350 0.835 91.350 4.280 ;
        RECT 92.190 0.835 92.730 4.280 ;
        RECT 93.570 0.835 94.570 4.280 ;
        RECT 95.410 0.835 95.950 4.280 ;
        RECT 96.790 0.835 97.790 4.280 ;
        RECT 98.630 0.835 99.170 4.280 ;
        RECT 100.010 0.835 101.010 4.280 ;
        RECT 101.850 0.835 102.390 4.280 ;
        RECT 103.230 0.835 104.230 4.280 ;
        RECT 105.070 0.835 105.610 4.280 ;
        RECT 106.450 0.835 107.450 4.280 ;
        RECT 108.290 0.835 108.830 4.280 ;
        RECT 109.670 0.835 110.670 4.280 ;
        RECT 111.510 0.835 112.050 4.280 ;
        RECT 112.890 0.835 113.890 4.280 ;
        RECT 114.730 0.835 115.270 4.280 ;
        RECT 116.110 0.835 117.110 4.280 ;
        RECT 117.950 0.835 118.490 4.280 ;
        RECT 119.330 0.835 120.330 4.280 ;
        RECT 121.170 0.835 121.710 4.280 ;
        RECT 122.550 0.835 123.090 4.280 ;
        RECT 123.930 0.835 124.930 4.280 ;
        RECT 125.770 0.835 126.310 4.280 ;
        RECT 127.150 0.835 128.150 4.280 ;
        RECT 128.990 0.835 129.530 4.280 ;
        RECT 130.370 0.835 131.370 4.280 ;
        RECT 132.210 0.835 132.750 4.280 ;
        RECT 133.590 0.835 134.590 4.280 ;
        RECT 135.430 0.835 135.970 4.280 ;
        RECT 136.810 0.835 137.810 4.280 ;
        RECT 138.650 0.835 139.190 4.280 ;
        RECT 140.030 0.835 141.030 4.280 ;
        RECT 141.870 0.835 142.410 4.280 ;
        RECT 143.250 0.835 144.250 4.280 ;
        RECT 145.090 0.835 145.630 4.280 ;
        RECT 146.470 0.835 147.470 4.280 ;
        RECT 148.310 0.835 148.850 4.280 ;
        RECT 149.690 0.835 150.690 4.280 ;
        RECT 151.530 0.835 152.070 4.280 ;
        RECT 152.910 0.835 153.910 4.280 ;
        RECT 154.750 0.835 155.290 4.280 ;
        RECT 156.130 0.835 157.130 4.280 ;
        RECT 157.970 0.835 158.510 4.280 ;
        RECT 159.350 0.835 160.350 4.280 ;
        RECT 161.190 0.835 161.730 4.280 ;
        RECT 162.570 0.835 163.110 4.280 ;
        RECT 163.950 0.835 164.950 4.280 ;
        RECT 165.790 0.835 166.330 4.280 ;
        RECT 167.170 0.835 168.170 4.280 ;
        RECT 169.010 0.835 169.550 4.280 ;
        RECT 170.390 0.835 171.390 4.280 ;
        RECT 172.230 0.835 172.770 4.280 ;
        RECT 173.610 0.835 174.610 4.280 ;
        RECT 175.450 0.835 175.990 4.280 ;
        RECT 176.830 0.835 177.830 4.280 ;
        RECT 178.670 0.835 179.210 4.280 ;
        RECT 180.050 0.835 181.050 4.280 ;
        RECT 181.890 0.835 182.430 4.280 ;
        RECT 183.270 0.835 184.270 4.280 ;
        RECT 185.110 0.835 185.650 4.280 ;
        RECT 186.490 0.835 187.490 4.280 ;
        RECT 188.330 0.835 188.870 4.280 ;
        RECT 189.710 0.835 190.710 4.280 ;
        RECT 191.550 0.835 192.090 4.280 ;
        RECT 192.930 0.835 193.930 4.280 ;
        RECT 194.770 0.835 195.310 4.280 ;
        RECT 196.150 0.835 197.150 4.280 ;
        RECT 197.990 0.835 198.530 4.280 ;
        RECT 199.370 0.835 200.370 4.280 ;
        RECT 201.210 0.835 201.750 4.280 ;
        RECT 202.590 0.835 203.130 4.280 ;
        RECT 203.970 0.835 204.970 4.280 ;
        RECT 205.810 0.835 206.350 4.280 ;
        RECT 207.190 0.835 208.190 4.280 ;
        RECT 209.030 0.835 209.570 4.280 ;
        RECT 210.410 0.835 211.410 4.280 ;
        RECT 212.250 0.835 212.790 4.280 ;
        RECT 213.630 0.835 214.630 4.280 ;
        RECT 215.470 0.835 216.010 4.280 ;
        RECT 216.850 0.835 217.850 4.280 ;
        RECT 218.690 0.835 219.230 4.280 ;
        RECT 220.070 0.835 221.070 4.280 ;
        RECT 221.910 0.835 222.450 4.280 ;
        RECT 223.290 0.835 224.290 4.280 ;
        RECT 225.130 0.835 225.670 4.280 ;
        RECT 226.510 0.835 227.510 4.280 ;
        RECT 228.350 0.835 228.890 4.280 ;
        RECT 229.730 0.835 230.730 4.280 ;
        RECT 231.570 0.835 232.110 4.280 ;
        RECT 232.950 0.835 233.950 4.280 ;
        RECT 234.790 0.835 235.330 4.280 ;
        RECT 236.170 0.835 237.170 4.280 ;
        RECT 238.010 0.835 238.550 4.280 ;
        RECT 239.390 0.835 240.390 4.280 ;
        RECT 241.230 0.835 241.770 4.280 ;
        RECT 242.610 0.835 243.150 4.280 ;
        RECT 243.990 0.835 244.990 4.280 ;
        RECT 245.830 0.835 246.370 4.280 ;
        RECT 247.210 0.835 248.210 4.280 ;
        RECT 249.050 0.835 249.590 4.280 ;
        RECT 250.430 0.835 251.430 4.280 ;
        RECT 252.270 0.835 252.810 4.280 ;
        RECT 253.650 0.835 254.650 4.280 ;
        RECT 255.490 0.835 256.030 4.280 ;
        RECT 256.870 0.835 257.870 4.280 ;
        RECT 258.710 0.835 259.250 4.280 ;
        RECT 260.090 0.835 261.090 4.280 ;
        RECT 261.930 0.835 262.470 4.280 ;
        RECT 263.310 0.835 264.310 4.280 ;
        RECT 265.150 0.835 265.690 4.280 ;
        RECT 266.530 0.835 267.530 4.280 ;
        RECT 268.370 0.835 268.910 4.280 ;
        RECT 269.750 0.835 270.750 4.280 ;
        RECT 271.590 0.835 272.130 4.280 ;
        RECT 272.970 0.835 273.970 4.280 ;
        RECT 274.810 0.835 275.350 4.280 ;
        RECT 276.190 0.835 277.190 4.280 ;
        RECT 278.030 0.835 278.570 4.280 ;
        RECT 279.410 0.835 280.410 4.280 ;
        RECT 281.250 0.835 281.790 4.280 ;
        RECT 282.630 0.835 283.170 4.280 ;
        RECT 284.010 0.835 285.010 4.280 ;
        RECT 285.850 0.835 286.390 4.280 ;
        RECT 287.230 0.835 288.230 4.280 ;
        RECT 289.070 0.835 289.610 4.280 ;
        RECT 290.450 0.835 291.450 4.280 ;
        RECT 292.290 0.835 292.830 4.280 ;
        RECT 293.670 0.835 294.670 4.280 ;
        RECT 295.510 0.835 296.050 4.280 ;
        RECT 296.890 0.835 297.890 4.280 ;
        RECT 298.730 0.835 299.270 4.280 ;
        RECT 300.110 0.835 301.110 4.280 ;
        RECT 301.950 0.835 302.490 4.280 ;
        RECT 303.330 0.835 304.330 4.280 ;
        RECT 305.170 0.835 305.710 4.280 ;
        RECT 306.550 0.835 307.550 4.280 ;
        RECT 308.390 0.835 308.930 4.280 ;
        RECT 309.770 0.835 310.770 4.280 ;
        RECT 311.610 0.835 312.150 4.280 ;
        RECT 312.990 0.835 313.990 4.280 ;
        RECT 314.830 0.835 315.370 4.280 ;
        RECT 316.210 0.835 317.210 4.280 ;
        RECT 318.050 0.835 318.590 4.280 ;
        RECT 319.430 0.835 320.430 4.280 ;
        RECT 321.270 0.835 321.810 4.280 ;
        RECT 322.650 0.835 323.190 4.280 ;
        RECT 324.030 0.835 325.030 4.280 ;
        RECT 325.870 0.835 326.410 4.280 ;
        RECT 327.250 0.835 328.250 4.280 ;
        RECT 329.090 0.835 329.630 4.280 ;
        RECT 330.470 0.835 331.470 4.280 ;
        RECT 332.310 0.835 332.850 4.280 ;
        RECT 333.690 0.835 334.690 4.280 ;
        RECT 335.530 0.835 336.070 4.280 ;
        RECT 336.910 0.835 337.910 4.280 ;
        RECT 338.750 0.835 339.290 4.280 ;
        RECT 340.130 0.835 341.130 4.280 ;
        RECT 341.970 0.835 342.510 4.280 ;
        RECT 343.350 0.835 344.350 4.280 ;
        RECT 345.190 0.835 345.730 4.280 ;
        RECT 346.570 0.835 347.570 4.280 ;
        RECT 348.410 0.835 348.950 4.280 ;
        RECT 349.790 0.835 350.790 4.280 ;
        RECT 351.630 0.835 352.170 4.280 ;
        RECT 353.010 0.835 354.010 4.280 ;
        RECT 354.850 0.835 355.390 4.280 ;
        RECT 356.230 0.835 357.230 4.280 ;
        RECT 358.070 0.835 358.610 4.280 ;
        RECT 359.450 0.835 360.450 4.280 ;
        RECT 361.290 0.835 361.830 4.280 ;
        RECT 362.670 0.835 363.210 4.280 ;
        RECT 364.050 0.835 365.050 4.280 ;
        RECT 365.890 0.835 366.430 4.280 ;
        RECT 367.270 0.835 368.270 4.280 ;
        RECT 369.110 0.835 369.650 4.280 ;
        RECT 370.490 0.835 371.490 4.280 ;
        RECT 372.330 0.835 372.870 4.280 ;
        RECT 373.710 0.835 374.710 4.280 ;
        RECT 375.550 0.835 376.090 4.280 ;
        RECT 376.930 0.835 377.930 4.280 ;
        RECT 378.770 0.835 379.310 4.280 ;
        RECT 380.150 0.835 381.150 4.280 ;
        RECT 381.990 0.835 382.530 4.280 ;
        RECT 383.370 0.835 384.370 4.280 ;
        RECT 385.210 0.835 385.750 4.280 ;
        RECT 386.590 0.835 387.590 4.280 ;
        RECT 388.430 0.835 388.970 4.280 ;
        RECT 389.810 0.835 390.810 4.280 ;
        RECT 391.650 0.835 392.190 4.280 ;
        RECT 393.030 0.835 394.030 4.280 ;
        RECT 394.870 0.835 395.410 4.280 ;
        RECT 396.250 0.835 397.250 4.280 ;
        RECT 398.090 0.835 398.630 4.280 ;
      LAYER met3 ;
        RECT 4.400 398.120 395.600 398.985 ;
        RECT 4.400 397.480 396.000 398.120 ;
        RECT 4.400 396.760 395.600 397.480 ;
        RECT 4.000 396.120 395.600 396.760 ;
        RECT 4.400 396.080 395.600 396.120 ;
        RECT 4.400 395.440 396.000 396.080 ;
        RECT 4.400 393.360 395.600 395.440 ;
        RECT 4.000 392.720 395.600 393.360 ;
        RECT 4.400 392.680 395.600 392.720 ;
        RECT 4.400 392.040 396.000 392.680 ;
        RECT 4.400 390.640 395.600 392.040 ;
        RECT 4.400 390.000 396.000 390.640 ;
        RECT 4.400 389.960 395.600 390.000 ;
        RECT 4.000 389.320 395.600 389.960 ;
        RECT 4.400 387.240 395.600 389.320 ;
        RECT 4.400 386.600 396.000 387.240 ;
        RECT 4.400 386.560 395.600 386.600 ;
        RECT 4.000 385.920 395.600 386.560 ;
        RECT 4.400 385.200 395.600 385.920 ;
        RECT 4.400 384.560 396.000 385.200 ;
        RECT 4.400 383.160 395.600 384.560 ;
        RECT 4.000 382.520 396.000 383.160 ;
        RECT 4.400 379.760 395.600 382.520 ;
        RECT 4.000 379.120 396.000 379.760 ;
        RECT 4.400 377.720 395.600 379.120 ;
        RECT 4.400 377.080 396.000 377.720 ;
        RECT 4.400 376.360 395.600 377.080 ;
        RECT 4.000 375.720 395.600 376.360 ;
        RECT 4.400 374.320 395.600 375.720 ;
        RECT 4.400 373.680 396.000 374.320 ;
        RECT 4.400 372.960 395.600 373.680 ;
        RECT 4.000 372.320 395.600 372.960 ;
        RECT 4.400 372.280 395.600 372.320 ;
        RECT 4.400 371.640 396.000 372.280 ;
        RECT 4.400 370.240 395.600 371.640 ;
        RECT 4.400 369.600 396.000 370.240 ;
        RECT 4.400 369.560 395.600 369.600 ;
        RECT 4.000 368.920 395.600 369.560 ;
        RECT 4.400 366.840 395.600 368.920 ;
        RECT 4.400 366.200 396.000 366.840 ;
        RECT 4.400 366.160 395.600 366.200 ;
        RECT 4.000 365.520 395.600 366.160 ;
        RECT 4.400 364.800 395.600 365.520 ;
        RECT 4.400 364.160 396.000 364.800 ;
        RECT 4.400 362.760 395.600 364.160 ;
        RECT 4.000 362.120 395.600 362.760 ;
        RECT 4.400 361.400 395.600 362.120 ;
        RECT 4.400 360.760 396.000 361.400 ;
        RECT 4.400 359.360 395.600 360.760 ;
        RECT 4.000 358.720 396.000 359.360 ;
        RECT 4.400 357.320 395.600 358.720 ;
        RECT 4.400 356.680 396.000 357.320 ;
        RECT 4.400 355.960 395.600 356.680 ;
        RECT 4.000 355.320 395.600 355.960 ;
        RECT 4.400 353.920 395.600 355.320 ;
        RECT 4.400 353.280 396.000 353.920 ;
        RECT 4.400 352.560 395.600 353.280 ;
        RECT 4.000 351.920 395.600 352.560 ;
        RECT 4.400 351.880 395.600 351.920 ;
        RECT 4.400 351.240 396.000 351.880 ;
        RECT 4.400 349.160 395.600 351.240 ;
        RECT 4.000 348.520 395.600 349.160 ;
        RECT 4.400 348.480 395.600 348.520 ;
        RECT 4.400 347.840 396.000 348.480 ;
        RECT 4.400 346.440 395.600 347.840 ;
        RECT 4.400 345.800 396.000 346.440 ;
        RECT 4.400 345.760 395.600 345.800 ;
        RECT 4.000 345.120 395.600 345.760 ;
        RECT 4.400 343.040 395.600 345.120 ;
        RECT 4.400 342.400 396.000 343.040 ;
        RECT 4.400 342.360 395.600 342.400 ;
        RECT 4.000 341.720 395.600 342.360 ;
        RECT 4.400 341.000 395.600 341.720 ;
        RECT 4.400 340.360 396.000 341.000 ;
        RECT 4.400 338.960 395.600 340.360 ;
        RECT 4.000 338.320 396.000 338.960 ;
        RECT 4.400 335.560 395.600 338.320 ;
        RECT 4.000 334.920 396.000 335.560 ;
        RECT 4.400 333.520 395.600 334.920 ;
        RECT 4.400 332.880 396.000 333.520 ;
        RECT 4.400 332.160 395.600 332.880 ;
        RECT 4.000 331.520 395.600 332.160 ;
        RECT 4.400 330.120 395.600 331.520 ;
        RECT 4.400 329.480 396.000 330.120 ;
        RECT 4.400 328.760 395.600 329.480 ;
        RECT 4.000 328.120 395.600 328.760 ;
        RECT 4.400 328.080 395.600 328.120 ;
        RECT 4.400 327.440 396.000 328.080 ;
        RECT 4.400 326.040 395.600 327.440 ;
        RECT 4.400 325.400 396.000 326.040 ;
        RECT 4.400 325.360 395.600 325.400 ;
        RECT 4.000 324.720 395.600 325.360 ;
        RECT 4.400 322.640 395.600 324.720 ;
        RECT 4.400 322.000 396.000 322.640 ;
        RECT 4.400 321.960 395.600 322.000 ;
        RECT 4.000 321.320 395.600 321.960 ;
        RECT 4.400 320.600 395.600 321.320 ;
        RECT 4.400 319.960 396.000 320.600 ;
        RECT 4.400 318.560 395.600 319.960 ;
        RECT 4.000 317.920 395.600 318.560 ;
        RECT 4.400 317.200 395.600 317.920 ;
        RECT 4.400 316.560 396.000 317.200 ;
        RECT 4.400 315.160 395.600 316.560 ;
        RECT 4.000 314.520 396.000 315.160 ;
        RECT 4.400 313.120 395.600 314.520 ;
        RECT 4.400 312.480 396.000 313.120 ;
        RECT 4.400 311.760 395.600 312.480 ;
        RECT 4.000 311.120 395.600 311.760 ;
        RECT 4.400 309.720 395.600 311.120 ;
        RECT 4.400 309.080 396.000 309.720 ;
        RECT 4.400 308.360 395.600 309.080 ;
        RECT 4.000 307.720 395.600 308.360 ;
        RECT 4.400 307.680 395.600 307.720 ;
        RECT 4.400 307.040 396.000 307.680 ;
        RECT 4.400 304.960 395.600 307.040 ;
        RECT 4.000 304.320 395.600 304.960 ;
        RECT 4.400 304.280 395.600 304.320 ;
        RECT 4.400 303.640 396.000 304.280 ;
        RECT 4.400 302.240 395.600 303.640 ;
        RECT 4.400 301.600 396.000 302.240 ;
        RECT 4.400 300.200 395.600 301.600 ;
        RECT 4.000 299.560 396.000 300.200 ;
        RECT 4.400 296.800 395.600 299.560 ;
        RECT 4.000 296.160 396.000 296.800 ;
        RECT 4.400 294.760 395.600 296.160 ;
        RECT 4.400 294.120 396.000 294.760 ;
        RECT 4.400 293.400 395.600 294.120 ;
        RECT 4.000 292.760 395.600 293.400 ;
        RECT 4.400 291.360 395.600 292.760 ;
        RECT 4.400 290.720 396.000 291.360 ;
        RECT 4.400 290.000 395.600 290.720 ;
        RECT 4.000 289.360 395.600 290.000 ;
        RECT 4.400 289.320 395.600 289.360 ;
        RECT 4.400 288.680 396.000 289.320 ;
        RECT 4.400 286.600 395.600 288.680 ;
        RECT 4.000 285.960 395.600 286.600 ;
        RECT 4.400 285.920 395.600 285.960 ;
        RECT 4.400 285.280 396.000 285.920 ;
        RECT 4.400 283.880 395.600 285.280 ;
        RECT 4.400 283.240 396.000 283.880 ;
        RECT 4.400 283.200 395.600 283.240 ;
        RECT 4.000 282.560 395.600 283.200 ;
        RECT 4.400 281.840 395.600 282.560 ;
        RECT 4.400 281.200 396.000 281.840 ;
        RECT 4.400 279.800 395.600 281.200 ;
        RECT 4.000 279.160 395.600 279.800 ;
        RECT 4.400 278.440 395.600 279.160 ;
        RECT 4.400 277.800 396.000 278.440 ;
        RECT 4.400 276.400 395.600 277.800 ;
        RECT 4.000 275.760 396.000 276.400 ;
        RECT 4.400 273.000 395.600 275.760 ;
        RECT 4.000 272.360 396.000 273.000 ;
        RECT 4.400 270.960 395.600 272.360 ;
        RECT 4.400 270.320 396.000 270.960 ;
        RECT 4.400 269.600 395.600 270.320 ;
        RECT 4.000 268.960 395.600 269.600 ;
        RECT 4.400 268.920 395.600 268.960 ;
        RECT 4.400 268.280 396.000 268.920 ;
        RECT 4.400 266.200 395.600 268.280 ;
        RECT 4.000 265.560 395.600 266.200 ;
        RECT 4.400 265.520 395.600 265.560 ;
        RECT 4.400 264.880 396.000 265.520 ;
        RECT 4.400 263.480 395.600 264.880 ;
        RECT 4.400 262.840 396.000 263.480 ;
        RECT 4.400 262.800 395.600 262.840 ;
        RECT 4.000 262.160 395.600 262.800 ;
        RECT 4.400 260.080 395.600 262.160 ;
        RECT 4.400 259.440 396.000 260.080 ;
        RECT 4.400 259.400 395.600 259.440 ;
        RECT 4.000 258.760 395.600 259.400 ;
        RECT 4.400 258.040 395.600 258.760 ;
        RECT 4.400 257.400 396.000 258.040 ;
        RECT 4.400 256.000 395.600 257.400 ;
        RECT 4.000 255.360 396.000 256.000 ;
        RECT 4.400 252.600 395.600 255.360 ;
        RECT 4.000 251.960 396.000 252.600 ;
        RECT 4.400 250.560 395.600 251.960 ;
        RECT 4.400 249.920 396.000 250.560 ;
        RECT 4.400 249.200 395.600 249.920 ;
        RECT 4.000 248.560 395.600 249.200 ;
        RECT 4.400 247.160 395.600 248.560 ;
        RECT 4.400 246.520 396.000 247.160 ;
        RECT 4.400 245.800 395.600 246.520 ;
        RECT 4.000 245.160 395.600 245.800 ;
        RECT 4.400 245.120 395.600 245.160 ;
        RECT 4.400 244.480 396.000 245.120 ;
        RECT 4.400 243.080 395.600 244.480 ;
        RECT 4.400 242.440 396.000 243.080 ;
        RECT 4.400 242.400 395.600 242.440 ;
        RECT 4.000 241.760 395.600 242.400 ;
        RECT 4.400 239.680 395.600 241.760 ;
        RECT 4.400 239.040 396.000 239.680 ;
        RECT 4.400 239.000 395.600 239.040 ;
        RECT 4.000 238.360 395.600 239.000 ;
        RECT 4.400 237.640 395.600 238.360 ;
        RECT 4.400 237.000 396.000 237.640 ;
        RECT 4.400 235.600 395.600 237.000 ;
        RECT 4.000 234.960 395.600 235.600 ;
        RECT 4.400 234.240 395.600 234.960 ;
        RECT 4.400 233.600 396.000 234.240 ;
        RECT 4.400 232.200 395.600 233.600 ;
        RECT 4.000 231.560 396.000 232.200 ;
        RECT 4.400 228.800 395.600 231.560 ;
        RECT 4.000 228.160 396.000 228.800 ;
        RECT 4.400 226.760 395.600 228.160 ;
        RECT 4.400 226.120 396.000 226.760 ;
        RECT 4.400 225.400 395.600 226.120 ;
        RECT 4.000 224.760 395.600 225.400 ;
        RECT 4.400 224.720 395.600 224.760 ;
        RECT 4.400 224.080 396.000 224.720 ;
        RECT 4.400 222.000 395.600 224.080 ;
        RECT 4.000 221.360 395.600 222.000 ;
        RECT 4.400 221.320 395.600 221.360 ;
        RECT 4.400 220.680 396.000 221.320 ;
        RECT 4.400 219.280 395.600 220.680 ;
        RECT 4.400 218.640 396.000 219.280 ;
        RECT 4.400 218.600 395.600 218.640 ;
        RECT 4.000 217.960 395.600 218.600 ;
        RECT 4.400 215.880 395.600 217.960 ;
        RECT 4.400 215.240 396.000 215.880 ;
        RECT 4.400 215.200 395.600 215.240 ;
        RECT 4.000 214.560 395.600 215.200 ;
        RECT 4.400 213.840 395.600 214.560 ;
        RECT 4.400 213.200 396.000 213.840 ;
        RECT 4.400 211.800 395.600 213.200 ;
        RECT 4.000 211.160 396.000 211.800 ;
        RECT 4.400 208.400 395.600 211.160 ;
        RECT 4.000 207.760 396.000 208.400 ;
        RECT 4.400 206.360 395.600 207.760 ;
        RECT 4.400 205.720 396.000 206.360 ;
        RECT 4.400 205.000 395.600 205.720 ;
        RECT 4.000 204.360 395.600 205.000 ;
        RECT 4.400 202.960 395.600 204.360 ;
        RECT 4.400 202.320 396.000 202.960 ;
        RECT 4.400 200.920 395.600 202.320 ;
        RECT 4.400 200.280 396.000 200.920 ;
        RECT 4.400 200.240 395.600 200.280 ;
        RECT 4.000 199.600 395.600 200.240 ;
        RECT 4.400 198.880 395.600 199.600 ;
        RECT 4.400 198.240 396.000 198.880 ;
        RECT 4.400 196.840 395.600 198.240 ;
        RECT 4.000 196.200 395.600 196.840 ;
        RECT 4.400 195.480 395.600 196.200 ;
        RECT 4.400 194.840 396.000 195.480 ;
        RECT 4.400 193.440 395.600 194.840 ;
        RECT 4.000 192.800 396.000 193.440 ;
        RECT 4.400 190.040 395.600 192.800 ;
        RECT 4.000 189.400 396.000 190.040 ;
        RECT 4.400 188.000 395.600 189.400 ;
        RECT 4.400 187.360 396.000 188.000 ;
        RECT 4.400 186.640 395.600 187.360 ;
        RECT 4.000 186.000 395.600 186.640 ;
        RECT 4.400 185.960 395.600 186.000 ;
        RECT 4.400 185.320 396.000 185.960 ;
        RECT 4.400 183.240 395.600 185.320 ;
        RECT 4.000 182.600 395.600 183.240 ;
        RECT 4.400 182.560 395.600 182.600 ;
        RECT 4.400 181.920 396.000 182.560 ;
        RECT 4.400 180.520 395.600 181.920 ;
        RECT 4.400 179.880 396.000 180.520 ;
        RECT 4.400 179.840 395.600 179.880 ;
        RECT 4.000 179.200 395.600 179.840 ;
        RECT 4.400 177.120 395.600 179.200 ;
        RECT 4.400 176.480 396.000 177.120 ;
        RECT 4.400 176.440 395.600 176.480 ;
        RECT 4.000 175.800 395.600 176.440 ;
        RECT 4.400 175.080 395.600 175.800 ;
        RECT 4.400 174.440 396.000 175.080 ;
        RECT 4.400 173.040 395.600 174.440 ;
        RECT 4.000 172.400 395.600 173.040 ;
        RECT 4.400 171.680 395.600 172.400 ;
        RECT 4.400 171.040 396.000 171.680 ;
        RECT 4.400 169.640 395.600 171.040 ;
        RECT 4.000 169.000 396.000 169.640 ;
        RECT 4.400 167.600 395.600 169.000 ;
        RECT 4.400 166.960 396.000 167.600 ;
        RECT 4.400 166.240 395.600 166.960 ;
        RECT 4.000 165.600 395.600 166.240 ;
        RECT 4.400 164.200 395.600 165.600 ;
        RECT 4.400 163.560 396.000 164.200 ;
        RECT 4.400 162.840 395.600 163.560 ;
        RECT 4.000 162.200 395.600 162.840 ;
        RECT 4.400 162.160 395.600 162.200 ;
        RECT 4.400 161.520 396.000 162.160 ;
        RECT 4.400 159.440 395.600 161.520 ;
        RECT 4.000 158.800 395.600 159.440 ;
        RECT 4.400 158.760 395.600 158.800 ;
        RECT 4.400 158.120 396.000 158.760 ;
        RECT 4.400 156.720 395.600 158.120 ;
        RECT 4.400 156.080 396.000 156.720 ;
        RECT 4.400 156.040 395.600 156.080 ;
        RECT 4.000 155.400 395.600 156.040 ;
        RECT 4.400 154.680 395.600 155.400 ;
        RECT 4.400 154.040 396.000 154.680 ;
        RECT 4.400 152.640 395.600 154.040 ;
        RECT 4.000 152.000 395.600 152.640 ;
        RECT 4.400 151.280 395.600 152.000 ;
        RECT 4.400 150.640 396.000 151.280 ;
        RECT 4.400 149.240 395.600 150.640 ;
        RECT 4.000 148.600 396.000 149.240 ;
        RECT 4.400 145.840 395.600 148.600 ;
        RECT 4.000 145.200 396.000 145.840 ;
        RECT 4.400 143.800 395.600 145.200 ;
        RECT 4.400 143.160 396.000 143.800 ;
        RECT 4.400 142.440 395.600 143.160 ;
        RECT 4.000 141.800 395.600 142.440 ;
        RECT 4.400 141.760 395.600 141.800 ;
        RECT 4.400 141.120 396.000 141.760 ;
        RECT 4.400 139.040 395.600 141.120 ;
        RECT 4.000 138.400 395.600 139.040 ;
        RECT 4.400 138.360 395.600 138.400 ;
        RECT 4.400 137.720 396.000 138.360 ;
        RECT 4.400 136.320 395.600 137.720 ;
        RECT 4.400 135.680 396.000 136.320 ;
        RECT 4.400 135.640 395.600 135.680 ;
        RECT 4.000 135.000 395.600 135.640 ;
        RECT 4.400 132.920 395.600 135.000 ;
        RECT 4.400 132.280 396.000 132.920 ;
        RECT 4.400 132.240 395.600 132.280 ;
        RECT 4.000 131.600 395.600 132.240 ;
        RECT 4.400 130.880 395.600 131.600 ;
        RECT 4.400 130.240 396.000 130.880 ;
        RECT 4.400 128.840 395.600 130.240 ;
        RECT 4.000 128.200 396.000 128.840 ;
        RECT 4.400 125.440 395.600 128.200 ;
        RECT 4.000 124.800 396.000 125.440 ;
        RECT 4.400 123.400 395.600 124.800 ;
        RECT 4.400 122.760 396.000 123.400 ;
        RECT 4.400 122.040 395.600 122.760 ;
        RECT 4.000 121.400 395.600 122.040 ;
        RECT 4.400 120.000 395.600 121.400 ;
        RECT 4.400 119.360 396.000 120.000 ;
        RECT 4.400 118.640 395.600 119.360 ;
        RECT 4.000 118.000 395.600 118.640 ;
        RECT 4.400 117.960 395.600 118.000 ;
        RECT 4.400 117.320 396.000 117.960 ;
        RECT 4.400 115.240 395.600 117.320 ;
        RECT 4.000 114.600 395.600 115.240 ;
        RECT 4.400 114.560 395.600 114.600 ;
        RECT 4.400 113.920 396.000 114.560 ;
        RECT 4.400 112.520 395.600 113.920 ;
        RECT 4.400 111.880 396.000 112.520 ;
        RECT 4.400 111.840 395.600 111.880 ;
        RECT 4.000 111.200 395.600 111.840 ;
        RECT 4.400 110.480 395.600 111.200 ;
        RECT 4.400 109.840 396.000 110.480 ;
        RECT 4.400 108.440 395.600 109.840 ;
        RECT 4.000 107.800 395.600 108.440 ;
        RECT 4.400 107.080 395.600 107.800 ;
        RECT 4.400 106.440 396.000 107.080 ;
        RECT 4.400 105.040 395.600 106.440 ;
        RECT 4.000 104.400 396.000 105.040 ;
        RECT 4.400 101.640 395.600 104.400 ;
        RECT 4.400 101.000 396.000 101.640 ;
        RECT 4.400 100.280 395.600 101.000 ;
        RECT 4.000 99.640 395.600 100.280 ;
        RECT 4.400 99.600 395.600 99.640 ;
        RECT 4.400 98.960 396.000 99.600 ;
        RECT 4.400 97.560 395.600 98.960 ;
        RECT 4.400 96.920 396.000 97.560 ;
        RECT 4.400 96.880 395.600 96.920 ;
        RECT 4.000 96.240 395.600 96.880 ;
        RECT 4.400 94.160 395.600 96.240 ;
        RECT 4.400 93.520 396.000 94.160 ;
        RECT 4.400 93.480 395.600 93.520 ;
        RECT 4.000 92.840 395.600 93.480 ;
        RECT 4.400 92.120 395.600 92.840 ;
        RECT 4.400 91.480 396.000 92.120 ;
        RECT 4.400 90.080 395.600 91.480 ;
        RECT 4.000 89.440 395.600 90.080 ;
        RECT 4.400 88.720 395.600 89.440 ;
        RECT 4.400 88.080 396.000 88.720 ;
        RECT 4.400 86.680 395.600 88.080 ;
        RECT 4.000 86.040 396.000 86.680 ;
        RECT 4.400 84.640 395.600 86.040 ;
        RECT 4.400 84.000 396.000 84.640 ;
        RECT 4.400 83.280 395.600 84.000 ;
        RECT 4.000 82.640 395.600 83.280 ;
        RECT 4.400 81.240 395.600 82.640 ;
        RECT 4.400 80.600 396.000 81.240 ;
        RECT 4.400 79.880 395.600 80.600 ;
        RECT 4.000 79.240 395.600 79.880 ;
        RECT 4.400 79.200 395.600 79.240 ;
        RECT 4.400 78.560 396.000 79.200 ;
        RECT 4.400 76.480 395.600 78.560 ;
        RECT 4.000 75.840 395.600 76.480 ;
        RECT 4.400 75.800 395.600 75.840 ;
        RECT 4.400 75.160 396.000 75.800 ;
        RECT 4.400 73.760 395.600 75.160 ;
        RECT 4.400 73.120 396.000 73.760 ;
        RECT 4.400 73.080 395.600 73.120 ;
        RECT 4.000 72.440 395.600 73.080 ;
        RECT 4.400 71.720 395.600 72.440 ;
        RECT 4.400 71.080 396.000 71.720 ;
        RECT 4.400 69.680 395.600 71.080 ;
        RECT 4.000 69.040 395.600 69.680 ;
        RECT 4.400 68.320 395.600 69.040 ;
        RECT 4.400 67.680 396.000 68.320 ;
        RECT 4.400 66.280 395.600 67.680 ;
        RECT 4.000 65.640 396.000 66.280 ;
        RECT 4.400 62.880 395.600 65.640 ;
        RECT 4.000 62.240 396.000 62.880 ;
        RECT 4.400 60.840 395.600 62.240 ;
        RECT 4.400 60.200 396.000 60.840 ;
        RECT 4.400 59.480 395.600 60.200 ;
        RECT 4.000 58.840 395.600 59.480 ;
        RECT 4.400 57.440 395.600 58.840 ;
        RECT 4.400 56.800 396.000 57.440 ;
        RECT 4.400 56.080 395.600 56.800 ;
        RECT 4.000 55.440 395.600 56.080 ;
        RECT 4.400 55.400 395.600 55.440 ;
        RECT 4.400 54.760 396.000 55.400 ;
        RECT 4.400 53.360 395.600 54.760 ;
        RECT 4.400 52.720 396.000 53.360 ;
        RECT 4.400 52.680 395.600 52.720 ;
        RECT 4.000 52.040 395.600 52.680 ;
        RECT 4.400 49.960 395.600 52.040 ;
        RECT 4.400 49.320 396.000 49.960 ;
        RECT 4.400 49.280 395.600 49.320 ;
        RECT 4.000 48.640 395.600 49.280 ;
        RECT 4.400 47.920 395.600 48.640 ;
        RECT 4.400 47.280 396.000 47.920 ;
        RECT 4.400 45.880 395.600 47.280 ;
        RECT 4.000 45.240 395.600 45.880 ;
        RECT 4.400 44.520 395.600 45.240 ;
        RECT 4.400 43.880 396.000 44.520 ;
        RECT 4.400 42.480 395.600 43.880 ;
        RECT 4.000 41.840 396.000 42.480 ;
        RECT 4.400 40.440 395.600 41.840 ;
        RECT 4.400 39.800 396.000 40.440 ;
        RECT 4.400 39.080 395.600 39.800 ;
        RECT 4.000 38.440 395.600 39.080 ;
        RECT 4.400 37.040 395.600 38.440 ;
        RECT 4.400 36.400 396.000 37.040 ;
        RECT 4.400 35.680 395.600 36.400 ;
        RECT 4.000 35.040 395.600 35.680 ;
        RECT 4.400 35.000 395.600 35.040 ;
        RECT 4.400 34.360 396.000 35.000 ;
        RECT 4.400 32.280 395.600 34.360 ;
        RECT 4.000 31.640 395.600 32.280 ;
        RECT 4.400 31.600 395.600 31.640 ;
        RECT 4.400 30.960 396.000 31.600 ;
        RECT 4.400 29.560 395.600 30.960 ;
        RECT 4.400 28.920 396.000 29.560 ;
        RECT 4.400 28.880 395.600 28.920 ;
        RECT 4.000 28.240 395.600 28.880 ;
        RECT 4.400 27.520 395.600 28.240 ;
        RECT 4.400 26.880 396.000 27.520 ;
        RECT 4.400 25.480 395.600 26.880 ;
        RECT 4.000 24.840 395.600 25.480 ;
        RECT 4.400 24.120 395.600 24.840 ;
        RECT 4.400 23.480 396.000 24.120 ;
        RECT 4.400 22.080 395.600 23.480 ;
        RECT 4.000 21.440 396.000 22.080 ;
        RECT 4.400 18.680 395.600 21.440 ;
        RECT 4.000 18.040 396.000 18.680 ;
        RECT 4.400 16.640 395.600 18.040 ;
        RECT 4.400 16.000 396.000 16.640 ;
        RECT 4.400 15.280 395.600 16.000 ;
        RECT 4.000 14.640 395.600 15.280 ;
        RECT 4.400 14.600 395.600 14.640 ;
        RECT 4.400 13.960 396.000 14.600 ;
        RECT 4.400 11.880 395.600 13.960 ;
        RECT 4.000 11.240 395.600 11.880 ;
        RECT 4.400 11.200 395.600 11.240 ;
        RECT 4.400 10.560 396.000 11.200 ;
        RECT 4.400 9.160 395.600 10.560 ;
        RECT 4.400 8.520 396.000 9.160 ;
        RECT 4.400 8.480 395.600 8.520 ;
        RECT 4.000 7.840 395.600 8.480 ;
        RECT 4.400 5.760 395.600 7.840 ;
        RECT 4.400 5.120 396.000 5.760 ;
        RECT 4.400 5.080 395.600 5.120 ;
        RECT 4.000 4.440 395.600 5.080 ;
        RECT 4.400 3.720 395.600 4.440 ;
        RECT 4.400 3.080 396.000 3.720 ;
        RECT 4.400 0.855 395.600 3.080 ;
      LAYER met4 ;
        RECT 17.775 12.415 20.640 267.065 ;
        RECT 23.040 12.415 97.440 267.065 ;
        RECT 99.840 12.415 174.240 267.065 ;
        RECT 176.640 12.415 251.040 267.065 ;
        RECT 253.440 12.415 292.265 267.065 ;
  END
END chip_controller
END LIBRARY

