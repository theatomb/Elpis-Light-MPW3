VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO io_output_arbiter
  CLASS BLOCK ;
  FOREIGN io_output_arbiter ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 75.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END clk
  PIN data_core0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 71.000 3.130 75.000 ;
    END
  END data_core0[0]
  PIN data_core0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END data_core0[10]
  PIN data_core0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 32.680 75.000 33.280 ;
    END
  END data_core0[11]
  PIN data_core0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 71.000 26.130 75.000 ;
    END
  END data_core0[12]
  PIN data_core0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END data_core0[13]
  PIN data_core0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END data_core0[14]
  PIN data_core0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 71.000 31.650 75.000 ;
    END
  END data_core0[15]
  PIN data_core0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END data_core0[16]
  PIN data_core0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END data_core0[17]
  PIN data_core0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END data_core0[18]
  PIN data_core0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 71.000 49.130 75.000 ;
    END
  END data_core0[19]
  PIN data_core0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END data_core0[1]
  PIN data_core0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END data_core0[20]
  PIN data_core0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END data_core0[21]
  PIN data_core0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END data_core0[22]
  PIN data_core0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END data_core0[23]
  PIN data_core0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 59.200 75.000 59.800 ;
    END
  END data_core0[24]
  PIN data_core0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 68.040 75.000 68.640 ;
    END
  END data_core0[25]
  PIN data_core0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 72.120 75.000 72.720 ;
    END
  END data_core0[26]
  PIN data_core0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END data_core0[27]
  PIN data_core0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END data_core0[28]
  PIN data_core0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END data_core0[29]
  PIN data_core0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 71.000 8.650 75.000 ;
    END
  END data_core0[2]
  PIN data_core0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END data_core0[30]
  PIN data_core0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END data_core0[31]
  PIN data_core0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 6.160 75.000 6.760 ;
    END
  END data_core0[3]
  PIN data_core0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 71.000 14.630 75.000 ;
    END
  END data_core0[4]
  PIN data_core0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END data_core0[5]
  PIN data_core0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END data_core0[6]
  PIN data_core0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 15.000 75.000 15.600 ;
    END
  END data_core0[7]
  PIN data_core0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END data_core0[8]
  PIN data_core0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 27.920 75.000 28.520 ;
    END
  END data_core0[9]
  PIN is_ready_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END is_ready_core0
  PIN print_hex_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END print_hex_enable
  PIN print_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END print_output[0]
  PIN print_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END print_output[10]
  PIN print_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 36.760 75.000 37.360 ;
    END
  END print_output[11]
  PIN print_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 41.520 75.000 42.120 ;
    END
  END print_output[12]
  PIN print_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END print_output[13]
  PIN print_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END print_output[14]
  PIN print_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 45.600 75.000 46.200 ;
    END
  END print_output[15]
  PIN print_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 71.000 37.630 75.000 ;
    END
  END print_output[16]
  PIN print_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 71.000 43.150 75.000 ;
    END
  END print_output[17]
  PIN print_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END print_output[18]
  PIN print_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 50.360 75.000 50.960 ;
    END
  END print_output[19]
  PIN print_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END print_output[1]
  PIN print_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END print_output[20]
  PIN print_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END print_output[21]
  PIN print_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END print_output[22]
  PIN print_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 54.440 75.000 55.040 ;
    END
  END print_output[23]
  PIN print_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 63.280 75.000 63.880 ;
    END
  END print_output[24]
  PIN print_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END print_output[25]
  PIN print_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END print_output[26]
  PIN print_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 71.000 54.650 75.000 ;
    END
  END print_output[27]
  PIN print_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 71.000 60.630 75.000 ;
    END
  END print_output[28]
  PIN print_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 71.000 66.150 75.000 ;
    END
  END print_output[29]
  PIN print_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 2.080 75.000 2.680 ;
    END
  END print_output[2]
  PIN print_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 71.000 72.130 75.000 ;
    END
  END print_output[30]
  PIN print_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END print_output[31]
  PIN print_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END print_output[3]
  PIN print_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 71.000 20.150 75.000 ;
    END
  END print_output[4]
  PIN print_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END print_output[5]
  PIN print_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 10.240 75.000 10.840 ;
    END
  END print_output[6]
  PIN print_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 19.080 75.000 19.680 ;
    END
  END print_output[7]
  PIN print_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 23.840 75.000 24.440 ;
    END
  END print_output[8]
  PIN print_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END print_output[9]
  PIN req_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END req_core0
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.380 10.640 16.980 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.700 10.640 38.300 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.020 10.640 59.620 62.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.040 10.640 27.640 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.360 10.640 48.960 62.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 2.465 71.155 68.255 ;
      LAYER met1 ;
        RECT 1.910 2.420 73.070 68.300 ;
      LAYER met2 ;
        RECT 1.940 70.720 2.570 72.605 ;
        RECT 3.410 70.720 8.090 72.605 ;
        RECT 8.930 70.720 14.070 72.605 ;
        RECT 14.910 70.720 19.590 72.605 ;
        RECT 20.430 70.720 25.570 72.605 ;
        RECT 26.410 70.720 31.090 72.605 ;
        RECT 31.930 70.720 37.070 72.605 ;
        RECT 37.910 70.720 42.590 72.605 ;
        RECT 43.430 70.720 48.570 72.605 ;
        RECT 49.410 70.720 54.090 72.605 ;
        RECT 54.930 70.720 60.070 72.605 ;
        RECT 60.910 70.720 65.590 72.605 ;
        RECT 66.430 70.720 71.570 72.605 ;
        RECT 72.410 70.720 73.040 72.605 ;
        RECT 1.940 4.280 73.040 70.720 ;
        RECT 2.490 1.515 5.330 4.280 ;
        RECT 6.170 1.515 9.470 4.280 ;
        RECT 10.310 1.515 13.150 4.280 ;
        RECT 13.990 1.515 17.290 4.280 ;
        RECT 18.130 1.515 20.970 4.280 ;
        RECT 21.810 1.515 25.110 4.280 ;
        RECT 25.950 1.515 29.250 4.280 ;
        RECT 30.090 1.515 32.930 4.280 ;
        RECT 33.770 1.515 37.070 4.280 ;
        RECT 37.910 1.515 40.750 4.280 ;
        RECT 41.590 1.515 44.890 4.280 ;
        RECT 45.730 1.515 48.570 4.280 ;
        RECT 49.410 1.515 52.710 4.280 ;
        RECT 53.550 1.515 56.850 4.280 ;
        RECT 57.690 1.515 60.530 4.280 ;
        RECT 61.370 1.515 64.670 4.280 ;
        RECT 65.510 1.515 68.350 4.280 ;
        RECT 69.190 1.515 72.490 4.280 ;
      LAYER met3 ;
        RECT 4.400 71.720 70.600 72.585 ;
        RECT 4.000 69.720 71.000 71.720 ;
        RECT 4.400 69.040 71.000 69.720 ;
        RECT 4.400 68.320 70.600 69.040 ;
        RECT 4.000 67.640 70.600 68.320 ;
        RECT 4.000 65.640 71.000 67.640 ;
        RECT 4.400 64.280 71.000 65.640 ;
        RECT 4.400 64.240 70.600 64.280 ;
        RECT 4.000 62.880 70.600 64.240 ;
        RECT 4.000 62.240 71.000 62.880 ;
        RECT 4.400 60.840 71.000 62.240 ;
        RECT 4.000 60.200 71.000 60.840 ;
        RECT 4.000 58.800 70.600 60.200 ;
        RECT 4.000 58.160 71.000 58.800 ;
        RECT 4.400 56.760 71.000 58.160 ;
        RECT 4.000 55.440 71.000 56.760 ;
        RECT 4.000 54.760 70.600 55.440 ;
        RECT 4.400 54.040 70.600 54.760 ;
        RECT 4.400 53.360 71.000 54.040 ;
        RECT 4.000 51.360 71.000 53.360 ;
        RECT 4.000 50.680 70.600 51.360 ;
        RECT 4.400 49.960 70.600 50.680 ;
        RECT 4.400 49.280 71.000 49.960 ;
        RECT 4.000 47.280 71.000 49.280 ;
        RECT 4.400 46.600 71.000 47.280 ;
        RECT 4.400 45.880 70.600 46.600 ;
        RECT 4.000 45.200 70.600 45.880 ;
        RECT 4.000 43.200 71.000 45.200 ;
        RECT 4.400 42.520 71.000 43.200 ;
        RECT 4.400 41.800 70.600 42.520 ;
        RECT 4.000 41.120 70.600 41.800 ;
        RECT 4.000 39.800 71.000 41.120 ;
        RECT 4.400 38.400 71.000 39.800 ;
        RECT 4.000 37.760 71.000 38.400 ;
        RECT 4.000 36.360 70.600 37.760 ;
        RECT 4.000 35.720 71.000 36.360 ;
        RECT 4.400 34.320 71.000 35.720 ;
        RECT 4.000 33.680 71.000 34.320 ;
        RECT 4.000 32.320 70.600 33.680 ;
        RECT 4.400 32.280 70.600 32.320 ;
        RECT 4.400 30.920 71.000 32.280 ;
        RECT 4.000 28.920 71.000 30.920 ;
        RECT 4.000 28.240 70.600 28.920 ;
        RECT 4.400 27.520 70.600 28.240 ;
        RECT 4.400 26.840 71.000 27.520 ;
        RECT 4.000 24.840 71.000 26.840 ;
        RECT 4.400 23.440 70.600 24.840 ;
        RECT 4.000 20.760 71.000 23.440 ;
        RECT 4.400 20.080 71.000 20.760 ;
        RECT 4.400 19.360 70.600 20.080 ;
        RECT 4.000 18.680 70.600 19.360 ;
        RECT 4.000 17.360 71.000 18.680 ;
        RECT 4.400 16.000 71.000 17.360 ;
        RECT 4.400 15.960 70.600 16.000 ;
        RECT 4.000 14.600 70.600 15.960 ;
        RECT 4.000 13.280 71.000 14.600 ;
        RECT 4.400 11.880 71.000 13.280 ;
        RECT 4.000 11.240 71.000 11.880 ;
        RECT 4.000 9.880 70.600 11.240 ;
        RECT 4.400 9.840 70.600 9.880 ;
        RECT 4.400 8.480 71.000 9.840 ;
        RECT 4.000 7.160 71.000 8.480 ;
        RECT 4.000 5.800 70.600 7.160 ;
        RECT 4.400 5.760 70.600 5.800 ;
        RECT 4.400 4.400 71.000 5.760 ;
        RECT 4.000 3.080 71.000 4.400 ;
        RECT 4.000 2.400 70.600 3.080 ;
        RECT 4.400 1.680 70.600 2.400 ;
        RECT 4.400 1.535 71.000 1.680 ;
  END
END io_output_arbiter
END LIBRARY

