* NGSPICE file created from storebuffer.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

.subckt storebuffer addr_in[0] addr_in[10] addr_in[11] addr_in[12] addr_in[13] addr_in[14]
+ addr_in[15] addr_in[16] addr_in[17] addr_in[18] addr_in[19] addr_in[1] addr_in[20]
+ addr_in[21] addr_in[22] addr_in[23] addr_in[24] addr_in[25] addr_in[26] addr_in[27]
+ addr_in[28] addr_in[29] addr_in[2] addr_in[30] addr_in[31] addr_in[3] addr_in[4]
+ addr_in[5] addr_in[6] addr_in[7] addr_in[8] addr_in[9] addr_out[0] addr_out[10]
+ addr_out[11] addr_out[12] addr_out[13] addr_out[14] addr_out[15] addr_out[16] addr_out[17]
+ addr_out[18] addr_out[19] addr_out[1] addr_out[20] addr_out[21] addr_out[22] addr_out[23]
+ addr_out[24] addr_out[25] addr_out[26] addr_out[27] addr_out[28] addr_out[29] addr_out[2]
+ addr_out[30] addr_out[31] addr_out[3] addr_out[4] addr_out[5] addr_out[6] addr_out[7]
+ addr_out[8] addr_out[9] clk data_in[0] data_in[10] data_in[11] data_in[12] data_in[13]
+ data_in[14] data_in[15] data_in[16] data_in[17] data_in[18] data_in[19] data_in[1]
+ data_in[20] data_in[21] data_in[22] data_in[23] data_in[24] data_in[25] data_in[26]
+ data_in[27] data_in[28] data_in[29] data_in[2] data_in[30] data_in[31] data_in[3]
+ data_in[4] data_in[5] data_in[6] data_in[7] data_in[8] data_in[9] data_out[0] data_out[10]
+ data_out[11] data_out[12] data_out[13] data_out[14] data_out[15] data_out[16] data_out[17]
+ data_out[18] data_out[19] data_out[1] data_out[20] data_out[21] data_out[22] data_out[23]
+ data_out[24] data_out[25] data_out[26] data_out[27] data_out[28] data_out[29] data_out[2]
+ data_out[30] data_out[31] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7]
+ data_out[8] data_out[9] drain_out empty_out full_out hit_dtlb is_byte is_byte_out
+ is_data_to_cache reset sb_hit sb_re sb_we stall_dcache vccd1 vssd1
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2479__B1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3155_ _3148_/A _3148_/B _3148_/Y vssd1 vssd1 vccd1 vccd1 _3156_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3086_ _3090_/B _3090_/D _3081_/B vssd1 vssd1 vccd1 vccd1 _3086_/X sky130_fd_sc_hd__a21bo_1
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2455__A _2455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ _3988_/A vssd1 vssd1 vccd1 vccd1 _3988_/X sky130_fd_sc_hd__clkbuf_1
X_2939_ _2939_/A _2944_/B vssd1 vssd1 vccd1 vccd1 _2939_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4609_ _4706_/CLK _4609_/D vssd1 vssd1 vccd1 vccd1 _4609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3346__D _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3911_ _4470_/Q _3906_/X _2532_/A _3909_/X vssd1 vssd1 vccd1 vccd1 _4470_/D sky130_fd_sc_hd__a22o_1
XFILLER_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3842_ _3842_/A vssd1 vssd1 vccd1 vccd1 _4500_/D sky130_fd_sc_hd__clkbuf_1
X_3773_ _4546_/Q _3771_/X _2505_/A _3772_/X vssd1 vssd1 vccd1 vccd1 _4546_/D sky130_fd_sc_hd__a22o_1
X_2724_ _3150_/A _2724_/B vssd1 vssd1 vccd1 vccd1 _2781_/A sky130_fd_sc_hd__nor2_1
X_2655_ _2655_/A _2655_/B vssd1 vssd1 vccd1 vccd1 _2768_/B sky130_fd_sc_hd__or2_1
X_2586_ _4626_/Q vssd1 vssd1 vccd1 vccd1 _2655_/A sky130_fd_sc_hd__inv_2
X_4325_ _4076_/X _4420_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4325_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4256_ _4255_/X input57/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4256_/X sky130_fd_sc_hd__mux2_2
X_4187_ _4116_/X _2494_/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4187_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3207_ _2779_/X _3157_/X _3154_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3208_/C sky130_fd_sc_hd__o211ai_1
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3138_ _3137_/A _3137_/B _3137_/Y vssd1 vssd1 vccd1 vccd1 _3138_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3069_ _3069_/A _3179_/A vssd1 vssd1 vccd1 vccd1 _3075_/C sky130_fd_sc_hd__or2_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3744__A _3751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_31_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3654__A _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ _2434_/C _2347_/X _2431_/X _2443_/D _2439_/X vssd1 vssd1 vccd1 vccd1 _2440_/X
+ sky130_fd_sc_hd__o221a_1
X_2371_ _2244_/Y _4576_/Q _2368_/Y _2369_/Y _2370_/X vssd1 vssd1 vccd1 vccd1 _2378_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_68_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4110_/A vssd1 vssd1 vccd1 vccd1 _4110_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4041_ _4041_/A vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2854__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3825_ _4260_/X _4506_/Q _3952_/S vssd1 vssd1 vccd1 vccd1 _3826_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3756_ _4557_/Q _3750_/X input9/X _3751_/X vssd1 vssd1 vccd1 vccd1 _4557_/D sky130_fd_sc_hd__a22o_1
X_2707_ _4366_/X _2700_/A _4363_/X _2705_/X _2706_/Y vssd1 vssd1 vccd1 vccd1 _2709_/C
+ sky130_fd_sc_hd__a221o_1
X_3687_ _4603_/Q _3680_/X _2543_/A _3683_/X vssd1 vssd1 vccd1 vccd1 _4603_/D sky130_fd_sc_hd__a22o_1
X_2638_ _2638_/A _2638_/B vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__and2_1
X_2569_ _4630_/Q vssd1 vssd1 vccd1 vccd1 _2721_/B sky130_fd_sc_hd__inv_2
XFILLER_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4308_ _4307_/X _4369_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4308_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4239_ _4238_/X _4377_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4239_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2845__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4334__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2376__A2 _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input55_A data_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_2_0_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4244__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3610_ _4272_/X _4651_/Q _3952_/S vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__mux2_1
X_4590_ _4634_/CLK _4590_/D vssd1 vssd1 vccd1 vccd1 _4590_/Q sky130_fd_sc_hd__dfxtp_1
X_3541_ _3541_/A vssd1 vssd1 vccd1 vccd1 _4681_/D sky130_fd_sc_hd__clkbuf_1
X_3472_ _4213_/X _4712_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3473_/A sky130_fd_sc_hd__mux2_1
X_2423_ _3204_/A vssd1 vssd1 vccd1 vccd1 _2426_/A sky130_fd_sc_hd__clkbuf_2
X_2354_ _2354_/A vssd1 vssd1 vccd1 vccd1 _2355_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2285_ _2288_/B vssd1 vssd1 vccd1 vccd1 _2285_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4024_ input1/X _4034_/B _4026_/C vssd1 vssd1 vccd1 vccd1 _4024_/Y sky130_fd_sc_hd__nor3_1
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3252__B1 _2505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3808_ _4520_/Q _3802_/X _4391_/X _3807_/X vssd1 vssd1 vccd1 vccd1 _4520_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4427__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3739_ _4570_/Q _3734_/X _2532_/A _3737_/X vssd1 vssd1 vccd1 vccd1 _4570_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4329__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3243__B1 _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3794__A1 _4530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4418__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4239__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2809__B1 _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2283__A _4603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2972_ _4453_/Q _2971_/Y _2968_/B vssd1 vssd1 vccd1 vccd1 _2973_/B sky130_fd_sc_hd__o21ai_1
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2588__A2 _2507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4711_ _4734_/CLK _4711_/D vssd1 vssd1 vccd1 vccd1 _4711_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4409__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4642_ _4642_/CLK _4642_/D vssd1 vssd1 vccd1 vccd1 _4642_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4573_ _4752_/CLK _4573_/D vssd1 vssd1 vccd1 vccd1 _4573_/Q sky130_fd_sc_hd__dfxtp_1
X_3524_ _4278_/X _4688_/Q _3530_/S vssd1 vssd1 vccd1 vccd1 _3525_/A sky130_fd_sc_hd__mux2_1
X_3455_ _3455_/A vssd1 vssd1 vccd1 vccd1 _4720_/D sky130_fd_sc_hd__clkbuf_1
X_2406_ _4359_/X _2357_/Y _2358_/X vssd1 vssd1 vccd1 vccd1 _2407_/C sky130_fd_sc_hd__a21bo_1
XFILLER_39_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3386_ _4266_/X _4752_/Q _3408_/S vssd1 vssd1 vccd1 vccd1 _3387_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2337_ _2336_/A _2336_/B _2336_/X vssd1 vssd1 vccd1 vccd1 _2337_/X sky130_fd_sc_hd__a21bo_1
XFILLER_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2268_ _2266_/X _2267_/X _2262_/X _2263_/Y vssd1 vssd1 vccd1 vccd1 _2268_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4007_ _4207_/X _4007_/B vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__and2_1
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2199_ _3287_/A vssd1 vssd1 vccd1 vccd1 _2202_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3289__A _3341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2579__A2 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3700__A1 _4594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3700__B2 _3697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3898__S _3900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input18_A addr_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4192__A1 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output86_A _4530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ input7/X _3060_/A input6/X _3148_/A vssd1 vssd1 vccd1 vccd1 _3240_/X sky130_fd_sc_hd__a22o_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3171_ _2377_/Y _3169_/Y _4194_/X _3170_/B _3170_/Y vssd1 vssd1 vccd1 vccd1 _3171_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2955_ _2340_/A _2942_/X _4210_/X _2945_/Y vssd1 vssd1 vccd1 vccd1 _2955_/X sky130_fd_sc_hd__o22a_1
X_2886_ _2532_/A _2923_/A _2883_/Y _2885_/X _2803_/X vssd1 vssd1 vccd1 vccd1 _2886_/X
+ sky130_fd_sc_hd__o221a_1
X_4625_ _4625_/CLK _4625_/D vssd1 vssd1 vccd1 vccd1 _4625_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3556__B _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4556_ _4556_/CLK _4556_/D vssd1 vssd1 vccd1 vccd1 _4556_/Q sky130_fd_sc_hd__dfxtp_2
X_3507_ _3816_/A vssd1 vssd1 vccd1 vccd1 _3788_/A sky130_fd_sc_hd__buf_2
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4487_ _4733_/CLK _4487_/D vssd1 vssd1 vccd1 vccd1 _4487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3572__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3438_ _4266_/X _4727_/Q _3442_/S vssd1 vssd1 vccd1 vccd1 _3439_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2497__A1 _2500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3974_/A _3972_/A _4006_/B vssd1 vssd1 vccd1 vccd1 _4007_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__3694__B1 _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2651__A _4700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4342__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3466__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput75 _4520_/Q vssd1 vssd1 vccd1 vccd1 addr_out[13] sky130_fd_sc_hd__buf_2
Xoutput97 _4511_/Q vssd1 vssd1 vccd1 vccd1 addr_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__2488__A1 _2507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 _4530_/Q vssd1 vssd1 vccd1 vccd1 addr_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3685__B1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output124_A _4502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3079__D _3119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2740_ _2651_/Y _2591_/Y _2738_/X vssd1 vssd1 vccd1 vccd1 _2741_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__4252__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2671_ _2266_/X _2665_/X _2666_/X _2790_/A vssd1 vssd1 vccd1 vccd1 _2690_/B sky130_fd_sc_hd__o211ai_1
X_4410_ _4754_/Q _4704_/Q _4671_/Q _4617_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4410_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4341_ _4166_/X _4155_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4341_/X sky130_fd_sc_hd__mux2_4
XANTENNA__2715__A2 _2702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4272_ _4271_/X input50/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4272_/X sky130_fd_sc_hd__mux2_1
X_3223_ _3163_/Y _3174_/X _3223_/C _3223_/D vssd1 vssd1 vccd1 vccd1 _3223_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__2479__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154_ _3154_/A _3154_/B vssd1 vssd1 vccd1 vccd1 _3154_/X sky130_fd_sc_hd__or2_1
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3085_ _4341_/X _3094_/A _4352_/X _3084_/Y vssd1 vssd1 vccd1 vccd1 _3115_/A sky130_fd_sc_hd__a22o_1
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3987_ _4200_/X _3995_/B vssd1 vssd1 vccd1 vccd1 _3988_/A sky130_fd_sc_hd__and2_1
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2938_ _2949_/B _2938_/B vssd1 vssd1 vccd1 vccd1 _2944_/B sky130_fd_sc_hd__or2_1
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2471__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2869_ _4131_/A _4450_/Q _2513_/A _4449_/Q _2837_/X vssd1 vssd1 vccd1 vccd1 _2869_/Y
+ sky130_fd_sc_hd__a221oi_2
X_4608_ _4706_/CLK _4608_/D vssd1 vssd1 vccd1 vccd1 _4608_/Q sky130_fd_sc_hd__dfxtp_1
X_4539_ _4746_/CLK _4539_/D vssd1 vssd1 vccd1 vccd1 _4539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4337__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3658__B1 _2500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4247__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3910_ _4471_/Q _3906_/X _2535_/A _3909_/X vssd1 vssd1 vccd1 vccd1 _4471_/D sky130_fd_sc_hd__a22o_1
XANTENNA__2633__B2 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3841_ _4302_/X _4500_/Q _3841_/S vssd1 vssd1 vccd1 vccd1 _3842_/A sky130_fd_sc_hd__mux2_1
X_3772_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2723_ _4633_/Q _2722_/Y _2702_/B vssd1 vssd1 vccd1 vccd1 _2724_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2654_ _2654_/A _2753_/A _2752_/B _2756_/B vssd1 vssd1 vccd1 vccd1 _2655_/B sky130_fd_sc_hd__or4_2
XFILLER_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2585_ _4625_/Q vssd1 vssd1 vccd1 vccd1 _2654_/A sky130_fd_sc_hd__clkinv_2
XFILLER_99_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4324_ _4323_/X _4372_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4324_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4011__A _4013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4255_ _4039_/Y input57/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4255_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3649__B1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4186_ _4122_/X _2508_/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4186_/X sky130_fd_sc_hd__mux2_1
X_3206_ _2426_/A _3204_/B _2417_/X _3199_/X vssd1 vssd1 vccd1 vccd1 _3209_/C sky130_fd_sc_hd__a22o_1
XANTENNA__2872__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3137_ _3137_/A _3137_/B vssd1 vssd1 vccd1 vccd1 _3137_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3068_ _4546_/Q vssd1 vssd1 vccd1 vccd1 _3179_/A sky130_fd_sc_hd__inv_2
XFILLER_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3297__A _4769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3812__B1 _4388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2370_ _4665_/Q _4575_/Q vssd1 vssd1 vccd1 vccd1 _2370_/X sky130_fd_sc_hd__or2_1
XFILLER_96_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4040_ _3969_/A _3284_/B _3969_/B vssd1 vssd1 vccd1 vccd1 _4041_/A sky130_fd_sc_hd__o21ba_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2854__A1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3824_ _4507_/Q _3788_/A _4378_/X _3303_/A vssd1 vssd1 vccd1 vccd1 _4507_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3755_ _4558_/Q _3750_/X _2464_/A _3751_/X vssd1 vssd1 vccd1 vccd1 _4558_/D sky130_fd_sc_hd__a22o_1
X_3686_ _4604_/Q _3680_/X _2803_/A _3683_/X vssd1 vssd1 vccd1 vccd1 _4604_/D sky130_fd_sc_hd__a22o_1
X_2706_ _2953_/A _2706_/B vssd1 vssd1 vccd1 vccd1 _2706_/Y sky130_fd_sc_hd__nor2_1
X_2637_ _2637_/A _2637_/B _2637_/C _2637_/D vssd1 vssd1 vccd1 vccd1 _2637_/X sky130_fd_sc_hd__or4_1
XANTENNA__2542__B1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2568_ _2612_/B _2616_/B _2612_/A vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2499_ _4118_/A vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4307_ _4096_/X _4369_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4307_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4238_ _4048_/X _4377_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4238_/X sky130_fd_sc_hd__mux2_1
X_4169_ _4169_/A vssd1 vssd1 vccd1 vccd1 _4169_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__2845__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4390__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3270__A1 _2536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4350__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input48_A data_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4381__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2256__D _2318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2834__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3540_ _4292_/X _4681_/Q _3548_/S vssd1 vssd1 vccd1 vccd1 _3541_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4260__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3471_ _3471_/A vssd1 vssd1 vccd1 vccd1 _4713_/D sky130_fd_sc_hd__clkbuf_1
X_2422_ _4360_/X vssd1 vssd1 vccd1 vccd1 _3204_/A sky130_fd_sc_hd__inv_2
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2353_ _3154_/A vssd1 vssd1 vccd1 vccd1 _2353_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3604__S _3606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2284_ _2284_/A _2293_/A _2293_/B vssd1 vssd1 vccd1 vccd1 _2288_/B sky130_fd_sc_hd__or3_1
XFILLER_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4023_ input1/X _4033_/B _4026_/C vssd1 vssd1 vccd1 vccd1 _4023_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4372__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3252__A1 _2498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3807_ _3814_/A vssd1 vssd1 vccd1 vccd1 _3807_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4427__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3738_ _4571_/Q _3734_/X _2535_/A _3737_/X vssd1 vssd1 vccd1 vccd1 _4571_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3669_ _4215_/X _4613_/Q _3730_/S vssd1 vssd1 vccd1 vccd1 _3670_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_45_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3514__S _3514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2818__B2 _4467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4345__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3243__A1 _2507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3794__A2 _3788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4418__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3424__S _3586_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2809__A1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4255__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2971_ _2971_/A _2971_/B vssd1 vssd1 vccd1 vccd1 _2971_/Y sky130_fd_sc_hd__nor2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4760_/CLK _4710_/D vssd1 vssd1 vccd1 vccd1 _4710_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4409__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4641_ _4644_/CLK _4641_/D vssd1 vssd1 vccd1 vccd1 _4641_/Q sky130_fd_sc_hd__dfxtp_2
X_4572_ _4760_/CLK _4572_/D vssd1 vssd1 vccd1 vccd1 _4572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3523_ _3523_/A vssd1 vssd1 vccd1 vccd1 _4689_/D sky130_fd_sc_hd__clkbuf_1
X_3454_ _4280_/X _4720_/Q _3458_/S vssd1 vssd1 vccd1 vccd1 _3455_/A sky130_fd_sc_hd__mux2_1
X_2405_ _2367_/Y _2385_/X _2443_/A _2403_/C _2404_/Y vssd1 vssd1 vccd1 vccd1 _2405_/X
+ sky130_fd_sc_hd__o32a_1
X_3385_ _3430_/S vssd1 vssd1 vccd1 vccd1 _3408_/S sky130_fd_sc_hd__buf_2
X_2336_ _2336_/A _2336_/B vssd1 vssd1 vccd1 vccd1 _2336_/X sky130_fd_sc_hd__or2_1
XFILLER_84_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2267_ _2273_/B _2273_/D _2258_/B vssd1 vssd1 vccd1 vccd1 _2267_/X sky130_fd_sc_hd__a21bo_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4750_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4006_ _4039_/B _4006_/B vssd1 vssd1 vccd1 vccd1 _4006_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2474__A _2474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2198_ _4765_/Q vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__inv_2
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3289__B _3342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_1_0_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3700__A2 _3696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3943__A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output79_A _4524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3170_ _4194_/X _3170_/B vssd1 vssd1 vccd1 vccd1 _3170_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2954_ _4366_/X _2947_/A _4363_/X _2952_/X _2953_/Y vssd1 vssd1 vccd1 vccd1 _2956_/C
+ sky130_fd_sc_hd__a221o_1
X_2885_ _2819_/A _2884_/X _2819_/D vssd1 vssd1 vccd1 vccd1 _2885_/X sky130_fd_sc_hd__o21ba_1
X_4624_ _4625_/CLK _4624_/D vssd1 vssd1 vccd1 vccd1 _4624_/Q sky130_fd_sc_hd__dfxtp_1
X_4555_ _4556_/CLK _4555_/D vssd1 vssd1 vccd1 vccd1 _4555_/Q sky130_fd_sc_hd__dfxtp_2
X_3506_ _3506_/A vssd1 vssd1 vccd1 vccd1 _3816_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4486_ _4719_/CLK _4486_/D vssd1 vssd1 vccd1 vccd1 _4486_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3572__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3437_ _3437_/A vssd1 vssd1 vccd1 vccd1 _4728_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3694__A1 _4598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3368_ _3368_/A vssd1 vssd1 vccd1 vccd1 _4006_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _4591_/Q _2318_/Y _2309_/B vssd1 vssd1 vccd1 vccd1 _2319_/Y sky130_fd_sc_hd__o21ai_1
X_3299_ _3299_/A _4337_/S vssd1 vssd1 vccd1 vccd1 _4195_/S sky130_fd_sc_hd__nor2_2
XFILLER_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput76 _4521_/Q vssd1 vssd1 vccd1 vccd1 addr_out[14] sky130_fd_sc_hd__buf_2
XFILLER_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput87 _4531_/Q vssd1 vssd1 vccd1 vccd1 addr_out[24] sky130_fd_sc_hd__buf_2
Xoutput98 _4512_/Q vssd1 vssd1 vccd1 vccd1 addr_out[5] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A addr_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2670_ _2916_/A _2670_/B vssd1 vssd1 vccd1 vccd1 _2790_/A sky130_fd_sc_hd__or2_1
XFILLER_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4340_ _4339_/X input38/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4340_/X sky130_fd_sc_hd__mux2_1
X_4271_ _4033_/Y input50/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4271_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3222_ _3216_/D _3146_/X _3213_/X _3225_/D _3221_/X vssd1 vssd1 vccd1 vccd1 _3222_/X
+ sky130_fd_sc_hd__o221a_1
X_3153_ _4553_/Q _3152_/Y _3148_/B vssd1 vssd1 vccd1 vccd1 _3154_/B sky130_fd_sc_hd__o21ai_1
XFILLER_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3084_ _3090_/A _3081_/B _3082_/B vssd1 vssd1 vccd1 vccd1 _3084_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3986_ _4034_/B _3994_/B vssd1 vssd1 vccd1 vccd1 _3986_/Y sky130_fd_sc_hd__nor2_1
X_2937_ _2937_/A _2937_/B _2937_/C _2937_/D vssd1 vssd1 vccd1 vccd1 _3032_/A sky130_fd_sc_hd__or4_4
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2868_ _2863_/X _2866_/X _2867_/X vssd1 vssd1 vccd1 vccd1 _2868_/X sky130_fd_sc_hd__a21bo_2
X_4607_ _4706_/CLK _4607_/D vssd1 vssd1 vccd1 vccd1 _4607_/Q sky130_fd_sc_hd__dfxtp_1
X_2799_ _2799_/A _2799_/B vssd1 vssd1 vccd1 vccd1 _2800_/B sky130_fd_sc_hd__or2_1
X_4538_ _4695_/CLK _4538_/D vssd1 vssd1 vccd1 vccd1 _4538_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4469_ _4571_/CLK _4469_/D vssd1 vssd1 vccd1 vccd1 _4469_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3758__A _3772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4353__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4101__B _4103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2633__A2 _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4263__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3840_ _3840_/A vssd1 vssd1 vccd1 vccd1 _4501_/D sky130_fd_sc_hd__clkbuf_1
X_3771_ _3771_/A vssd1 vssd1 vccd1 vccd1 _3771_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2722_ _2722_/A _2722_/B vssd1 vssd1 vccd1 vccd1 _2722_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2653_ _2653_/A _2735_/A _2735_/B vssd1 vssd1 vccd1 vccd1 _2756_/B sky130_fd_sc_hd__or3_2
X_2584_ _4633_/Q _4136_/A _4632_/Q _2484_/A _2583_/X vssd1 vssd1 vccd1 vccd1 _2589_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4323_ _4078_/X _4372_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4323_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4011__B _4032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4254_ _4253_/X _3985_/A _4354_/S vssd1 vssd1 vccd1 vccd1 _4254_/X sky130_fd_sc_hd__mux2_2
XANTENNA__3649__B2 _3648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4185_ _4769_/Q vssd1 vssd1 vccd1 vccd1 _4185_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3205_ _2409_/X _3201_/X _3210_/A _3204_/X vssd1 vssd1 vccd1 vccd1 _3209_/B sky130_fd_sc_hd__o211ai_1
XFILLER_82_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3136_ _4349_/X vssd1 vssd1 vccd1 vccd1 _3136_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3067_ _4547_/Q vssd1 vssd1 vccd1 vccd1 _3069_/A sky130_fd_sc_hd__inv_2
XFILLER_27_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3821__B2 _3303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3821__A1 _4510_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3297__B _3297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3969_ _3969_/A _3969_/B vssd1 vssd1 vccd1 vccd1 _3970_/A sky130_fd_sc_hd__or2_1
XFILLER_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3888__A1 _4479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4348__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3812__A1 _4517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2615__A2 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4258__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3803__A1 _4524_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3803__B2 _3800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3823_ _4508_/Q _3788_/A _4379_/X _3303_/A vssd1 vssd1 vccd1 vccd1 _4508_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3754_ _4559_/Q _3750_/X _2455_/A _3751_/X vssd1 vssd1 vccd1 vccd1 _4559_/D sky130_fd_sc_hd__a22o_1
X_3685_ _4605_/Q _3680_/X _2532_/A _3683_/X vssd1 vssd1 vccd1 vccd1 _4605_/D sky130_fd_sc_hd__a22o_1
X_2705_ _4637_/Q _2704_/Y _2697_/B vssd1 vssd1 vccd1 vccd1 _2705_/X sky130_fd_sc_hd__o21a_1
X_2636_ _2636_/A _2638_/A _2636_/C _2638_/B vssd1 vssd1 vccd1 vccd1 _2637_/D sky130_fd_sc_hd__or4b_1
XANTENNA__4022__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2542__A1 _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3334__A3 _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2567_ _4637_/Q _2457_/A _4636_/Q _2466_/A vssd1 vssd1 vccd1 vccd1 _2612_/A sky130_fd_sc_hd__o22a_1
X_2498_ _2498_/A vssd1 vssd1 vccd1 vccd1 _4118_/A sky130_fd_sc_hd__inv_2
X_4306_ _4305_/X _4428_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4306_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4237_ _4236_/X _4001_/A _4354_/S vssd1 vssd1 vccd1 vccd1 _4237_/X sky130_fd_sc_hd__mux2_2
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ _4168_/A vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4390__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3119_ _3119_/A _3119_/B vssd1 vssd1 vccd1 vccd1 _3132_/B sky130_fd_sc_hd__or2_1
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4099_ _4429_/X _4103_/B vssd1 vssd1 vccd1 vccd1 _4100_/A sky130_fd_sc_hd__and2_1
XFILLER_70_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3270__A2 _4571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3771__A _3771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4286__A1 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4381__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4210__A1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3470_ _4340_/X _4713_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3471_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3681__A _3717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2421_ _2409_/X _2410_/Y _2415_/Y _2428_/B vssd1 vssd1 vccd1 vccd1 _2427_/B sky130_fd_sc_hd__o211ai_1
XANTENNA__3721__B1 _2500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2352_ _4361_/X vssd1 vssd1 vccd1 vccd1 _3154_/A sky130_fd_sc_hd__inv_2
X_2283_ _4603_/Q vssd1 vssd1 vccd1 vccd1 _2293_/A sky130_fd_sc_hd__inv_2
XFILLER_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4022_ input1/X _4032_/B _4026_/C vssd1 vssd1 vccd1 vccd1 _4022_/Y sky130_fd_sc_hd__nor3_1
XFILLER_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4372__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2827__A2 _4456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3806_ _4521_/Q _3802_/X _4392_/X _3800_/X vssd1 vssd1 vccd1 vccd1 _4521_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4201__A1 _3981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3737_ _3751_/A vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3668_ _3668_/A vssd1 vssd1 vccd1 vccd1 _4614_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_opt_1_0_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2619_ _4641_/Q _4152_/A _2563_/Y _2617_/X _2618_/X vssd1 vssd1 vccd1 vccd1 _2619_/X
+ sky130_fd_sc_hd__o221a_1
X_3599_ _3599_/A vssd1 vssd1 vccd1 vccd1 _3601_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3307__A3 _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3712__B1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2515__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4268__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3779__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4361__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3951__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input60_A data_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4259__A1 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3440__S _3442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2970_ _3150_/A _2970_/B vssd1 vssd1 vccd1 vccd1 _3024_/A sky130_fd_sc_hd__nor2_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4640_ _4644_/CLK _4640_/D vssd1 vssd1 vccd1 vccd1 _4640_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4271__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4571_ _4571_/CLK _4571_/D vssd1 vssd1 vccd1 vccd1 _4571_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3942__B1 _2507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3522_ _4276_/X _4689_/Q _3530_/S vssd1 vssd1 vccd1 vccd1 _3523_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3453_ _3453_/A vssd1 vssd1 vccd1 vccd1 _4721_/D sky130_fd_sc_hd__clkbuf_1
X_2404_ _2393_/X _2403_/A _2397_/X _2403_/D vssd1 vssd1 vccd1 vccd1 _2404_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3384_ _3569_/A _3576_/B _3588_/C vssd1 vssd1 vccd1 vccd1 _3430_/S sky130_fd_sc_hd__or3_4
X_2335_ _2327_/X _2329_/Y _2345_/A vssd1 vssd1 vccd1 vccd1 _2344_/A sky130_fd_sc_hd__o21ai_1
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2266_ _2266_/A vssd1 vssd1 vccd1 vccd1 _2266_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4005_ _4005_/A vssd1 vssd1 vccd1 vccd1 _4039_/B sky130_fd_sc_hd__clkinv_2
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3289__C _3289_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4769_ _4769_/CLK _4769_/D vssd1 vssd1 vccd1 vccd1 _4769_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__3933__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4356__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3924__B1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3381__D _3381_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4266__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_44_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2953_ _2953_/A _2953_/B vssd1 vssd1 vccd1 vccd1 _2953_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2884_ _2819_/C _2884_/B vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__and2b_1
XFILLER_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4623_ _4623_/CLK _4623_/D vssd1 vssd1 vccd1 vccd1 _4623_/Q sky130_fd_sc_hd__dfxtp_2
X_4554_ _4556_/CLK _4554_/D vssd1 vssd1 vccd1 vccd1 _4554_/Q sky130_fd_sc_hd__dfxtp_1
X_3505_ _3505_/A vssd1 vssd1 vccd1 vccd1 _4696_/D sky130_fd_sc_hd__clkbuf_1
X_4485_ _4719_/CLK _4485_/D vssd1 vssd1 vccd1 vccd1 _4485_/Q sky130_fd_sc_hd__dfxtp_2
X_3436_ _4264_/X _4728_/Q _3442_/S vssd1 vssd1 vccd1 vccd1 _3437_/A sky130_fd_sc_hd__mux2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _3367_/A _3392_/A vssd1 vssd1 vccd1 vccd1 _3368_/A sky130_fd_sc_hd__or2_1
XFILLER_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2318_ _2318_/A vssd1 vssd1 vccd1 vccd1 _2318_/Y sky130_fd_sc_hd__inv_2
X_3298_ _3298_/A vssd1 vssd1 vccd1 vccd1 _4337_/S sky130_fd_sc_hd__buf_12
X_2249_ _2249_/A _2249_/B vssd1 vssd1 vccd1 vccd1 _2250_/B sky130_fd_sc_hd__or2_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput77 _4522_/Q vssd1 vssd1 vccd1 vccd1 addr_out[15] sky130_fd_sc_hd__buf_2
Xoutput88 _4532_/Q vssd1 vssd1 vccd1 vccd1 addr_out[25] sky130_fd_sc_hd__buf_2
Xoutput99 _4513_/Q vssd1 vssd1 vccd1 vccd1 addr_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input23_A addr_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4398__A0 _4638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4270_ _4269_/X input51/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4270_/X sky130_fd_sc_hd__mux2_2
XFILLER_97_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3221_ _3217_/Y _3218_/X _3115_/D _3114_/A _3220_/Y vssd1 vssd1 vccd1 vccd1 _3221_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3152_ _3152_/A _3152_/B vssd1 vssd1 vccd1 vccd1 _3152_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3083_ _3089_/B _3082_/B _3082_/Y vssd1 vssd1 vccd1 vccd1 _3094_/A sky130_fd_sc_hd__a21oi_1
XFILLER_54_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3985_ _3985_/A vssd1 vssd1 vccd1 vccd1 _4034_/B sky130_fd_sc_hd__clkinv_2
X_2936_ _2936_/A _2936_/B _2936_/C _2936_/D vssd1 vssd1 vccd1 vccd1 _2937_/D sky130_fd_sc_hd__or4_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4025__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2867_ _4119_/A _4446_/Q _4120_/A _4447_/Q vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__o22a_1
X_4606_ _4649_/CLK _4606_/D vssd1 vssd1 vccd1 vccd1 _4606_/Q sky130_fd_sc_hd__dfxtp_1
X_2798_ _2798_/A _2798_/B _2798_/C _2798_/D vssd1 vssd1 vccd1 vccd1 _2799_/B sky130_fd_sc_hd__nor4_1
X_4537_ _4695_/CLK _4537_/D vssd1 vssd1 vccd1 vccd1 _4537_/Q sky130_fd_sc_hd__dfxtp_4
X_4468_ _4571_/CLK _4468_/D vssd1 vssd1 vccd1 vccd1 _4468_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3419_ _3419_/A vssd1 vssd1 vccd1 vccd1 _4736_/D sky130_fd_sc_hd__clkbuf_1
X_4399_ _4639_/Q _4596_/Q _4561_/Q _4461_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4399_/X sky130_fd_sc_hd__mux4_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2627__B1 _4642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2866__B1 _2505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2572__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3770_ _4547_/Q _3764_/X _2507_/A _3765_/X vssd1 vssd1 vccd1 vccd1 _4547_/D sky130_fd_sc_hd__a22o_1
X_2721_ _2721_/A _2721_/B _2725_/B vssd1 vssd1 vccd1 vccd1 _2722_/B sky130_fd_sc_hd__or3_1
X_2652_ _4619_/Q _4618_/Q _2651_/Y vssd1 vssd1 vccd1 vccd1 _2735_/B sky130_fd_sc_hd__o21ai_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2583_ _2649_/A input7/X _2722_/A input6/X vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__a22o_1
X_4322_ _4321_/X _4421_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4322_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4253_ _3988_/X _3985_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__mux2_1
X_3204_ _3204_/A _3204_/B vssd1 vssd1 vccd1 vccd1 _3204_/X sky130_fd_sc_hd__or2_1
XANTENNA__3649__A2 _3647_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4184_ _4773_/Q _3308_/Y _3964_/Y _3308_/A _2212_/X vssd1 vssd1 vccd1 vccd1 _4773_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3135_ _2327_/X _3131_/X _3144_/A vssd1 vssd1 vccd1 vccd1 _3143_/A sky130_fd_sc_hd__o21ai_1
X_3066_ _4544_/Q vssd1 vssd1 vccd1 vccd1 _3182_/A sky130_fd_sc_hd__inv_2
XFILLER_82_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3821__A2 _3816_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3968_ _4768_/Q vssd1 vssd1 vccd1 vccd1 _3968_/Y sky130_fd_sc_hd__inv_2
X_2919_ _2916_/A _2916_/B _2277_/Y _2918_/Y vssd1 vssd1 vccd1 vccd1 _2937_/C sky130_fd_sc_hd__a22o_1
X_3899_ _3899_/A vssd1 vssd1 vccd1 vccd1 _4474_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3594__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2938__A _2949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4364__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3679__A _3717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3264__B1 _3259_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4274__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3803__A2 _3802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3822_ _4509_/Q _3788_/A _4380_/X _3303_/A vssd1 vssd1 vccd1 vccd1 _4509_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _4560_/Q _3750_/X _2452_/A _3751_/X vssd1 vssd1 vccd1 vccd1 _4560_/D sky130_fd_sc_hd__a22o_1
X_3684_ _4606_/Q _3680_/X _2535_/A _3683_/X vssd1 vssd1 vccd1 vccd1 _4606_/D sky130_fd_sc_hd__a22o_1
X_2704_ _2704_/A _2704_/B vssd1 vssd1 vccd1 vccd1 _2704_/Y sky130_fd_sc_hd__nor2_1
X_2635_ _2667_/B _2815_/A _2668_/A _2816_/A vssd1 vssd1 vccd1 vccd1 _2638_/B sky130_fd_sc_hd__o22a_1
XANTENNA__4022__B _4032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4305_ _4098_/X _4428_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4305_/X sky130_fd_sc_hd__mux2_1
X_2566_ _4636_/Q _4147_/A _4635_/Q _4146_/A vssd1 vssd1 vccd1 vccd1 _2616_/B sky130_fd_sc_hd__a22o_1
X_2497_ _2500_/A _2247_/A _2492_/A _2246_/A vssd1 vssd1 vccd1 vccd1 _2497_/X sky130_fd_sc_hd__o22a_1
XFILLER_87_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ _4004_/X _4001_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _4236_/X sky130_fd_sc_hd__mux2_1
X_4167_ _4154_/A _4154_/B _4155_/B vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__a21bo_1
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3118_ _3118_/A _3118_/B vssd1 vssd1 vccd1 vccd1 _3118_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4098_ _4098_/A vssd1 vssd1 vccd1 vccd1 _4098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2493__A _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3049_ _4561_/Q vssd1 vssd1 vccd1 vccd1 _3137_/A sky130_fd_sc_hd__inv_2
XFILLER_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4359__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3246__B1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4107__B _4109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3438__S _3442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2420_ _2417_/X _2419_/X _2412_/X _2414_/X vssd1 vssd1 vccd1 vccd1 _2428_/B sky130_fd_sc_hd__o22a_1
XFILLER_89_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2351_ _3150_/A _2351_/B vssd1 vssd1 vccd1 vccd1 _2407_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4269__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2282_ _4604_/Q vssd1 vssd1 vccd1 vccd1 _2284_/A sky130_fd_sc_hd__inv_2
X_4021_ _4029_/C vssd1 vssd1 vccd1 vccd1 _4026_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3805_ _4522_/Q _3802_/X _4393_/X _3800_/X vssd1 vssd1 vccd1 vccd1 _4522_/D sky130_fd_sc_hd__a22o_1
X_3736_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3751_/A sky130_fd_sc_hd__buf_4
X_3667_ _4217_/X _4614_/Q _3730_/S vssd1 vssd1 vccd1 vccd1 _3668_/A sky130_fd_sc_hd__mux2_1
X_2618_ _4641_/Q _2446_/A _4640_/Q _4151_/A vssd1 vssd1 vccd1 vccd1 _2618_/X sky130_fd_sc_hd__a211o_1
X_3598_ _4354_/X _4353_/X _3598_/C vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__or3_1
X_2549_ _2549_/A _2551_/A _2549_/C _2551_/B vssd1 vssd1 vccd1 vccd1 _2550_/D sky130_fd_sc_hd__or4b_1
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4219_ _4218_/X _4373_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4219_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3779__B2 _3751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2451__A1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3951__B2 _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A data_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4570_ _4571_/CLK _4570_/D vssd1 vssd1 vccd1 vccd1 _4570_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3942__A1 _4447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3521_ _3536_/S vssd1 vssd1 vccd1 vccd1 _3530_/S sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_3_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3452_ _4278_/X _4721_/Q _3458_/S vssd1 vssd1 vccd1 vccd1 _3453_/A sky130_fd_sc_hd__mux2_1
X_2403_ _2403_/A _2403_/B _2403_/C _2403_/D vssd1 vssd1 vccd1 vccd1 _2443_/A sky130_fd_sc_hd__or4_4
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3383_ _3974_/A _3972_/A _4039_/C _3352_/A vssd1 vssd1 vccd1 vccd1 _3588_/C sky130_fd_sc_hd__o211a_1
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2334_ _3134_/A _2334_/B vssd1 vssd1 vccd1 vccd1 _2345_/A sky130_fd_sc_hd__or2_1
XFILLER_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2265_ _4345_/X vssd1 vssd1 vccd1 vccd1 _2266_/A sky130_fd_sc_hd__inv_2
XANTENNA__3458__A0 _4284_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4004_ _4004_/A vssd1 vssd1 vccd1 vccd1 _4004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4028__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3630__B1 _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4768_ _4773_/CLK _4768_/D vssd1 vssd1 vccd1 vccd1 _4768_/Q sky130_fd_sc_hd__dfxtp_1
X_3719_ _4581_/Q _3717_/X _2505_/A _3718_/X vssd1 vssd1 vccd1 vccd1 _4581_/D sky130_fd_sc_hd__a22o_1
X_4699_ _4750_/CLK _4699_/D vssd1 vssd1 vccd1 vccd1 _4699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3621__B1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3688__B1 _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2952_ _4459_/Q _2951_/Y _2944_/B vssd1 vssd1 vccd1 vccd1 _2952_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4282__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2883_ _2883_/A vssd1 vssd1 vccd1 vccd1 _2883_/Y sky130_fd_sc_hd__inv_2
X_4622_ _4623_/CLK _4622_/D vssd1 vssd1 vccd1 vccd1 _4622_/Q sky130_fd_sc_hd__dfxtp_1
X_4553_ _4556_/CLK _4553_/D vssd1 vssd1 vccd1 vccd1 _4553_/Q sky130_fd_sc_hd__dfxtp_1
X_4484_ _4733_/CLK _4484_/D vssd1 vssd1 vccd1 vccd1 _4484_/Q sky130_fd_sc_hd__dfxtp_1
X_3504_ _4264_/X _4696_/Q _3514_/S vssd1 vssd1 vccd1 vccd1 _3505_/A sky130_fd_sc_hd__mux2_1
X_3435_ _3435_/A vssd1 vssd1 vccd1 vccd1 _4729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4340__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3366_ input1/X _3366_/B vssd1 vssd1 vccd1 vccd1 _3392_/A sky130_fd_sc_hd__or2_1
XFILLER_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2317_/A vssd1 vssd1 vccd1 vccd1 _2317_/X sky130_fd_sc_hd__clkbuf_2
X_3297_ _4769_/Q _3297_/B vssd1 vssd1 vccd1 vccd1 _3298_/A sky130_fd_sc_hd__and2_1
X_2248_ _2248_/A _2248_/B vssd1 vssd1 vccd1 vccd1 _2249_/B sky130_fd_sc_hd__or2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4192__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput78 _4523_/Q vssd1 vssd1 vccd1 vccd1 addr_out[16] sky130_fd_sc_hd__buf_2
Xoutput89 _4533_/Q vssd1 vssd1 vccd1 vccd1 addr_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4367__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input16_A addr_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4398__A1 _4595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3300__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3220_ _3219_/Y _3111_/A _3114_/B _3114_/D vssd1 vssd1 vccd1 vccd1 _3220_/Y sky130_fd_sc_hd__a31oi_1
XANTENNA__3125__A2 _3119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3151_ _3151_/A vssd1 vssd1 vccd1 vccd1 _3152_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4277__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3082_ _3089_/B _3082_/B vssd1 vssd1 vccd1 vccd1 _3082_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ _3984_/A vssd1 vssd1 vccd1 vccd1 _3984_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2935_ _2925_/A _2925_/B _2301_/A _2932_/B vssd1 vssd1 vccd1 vccd1 _2936_/D sky130_fd_sc_hd__a22o_1
X_2866_ _2498_/A _2994_/A _2505_/A _2995_/A vssd1 vssd1 vccd1 vccd1 _2866_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4605_ _4649_/CLK _4605_/D vssd1 vssd1 vccd1 vccd1 _4605_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2797_ _2377_/A _2741_/A _2743_/X _2796_/X vssd1 vssd1 vccd1 vccd1 _2798_/B sky130_fd_sc_hd__o211ai_2
XFILLER_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4536_ _4649_/CLK _4536_/D vssd1 vssd1 vccd1 vccd1 _4536_/Q sky130_fd_sc_hd__dfxtp_1
X_4467_ _4571_/CLK _4467_/D vssd1 vssd1 vccd1 vccd1 _4467_/Q sky130_fd_sc_hd__dfxtp_2
X_4398_ _4638_/Q _4595_/Q _4560_/Q _4460_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4398_/X sky130_fd_sc_hd__mux4_1
X_3418_ _4290_/X _4736_/Q _3418_/S vssd1 vssd1 vccd1 vccd1 _3419_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input8_A addr_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4187__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3349_ _4367_/S _3349_/B vssd1 vssd1 vccd1 vccd1 _4339_/S sky130_fd_sc_hd__nor2_8
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2627__B2 _4153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_43_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2866__A1 _2498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output122_A _4500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3815__B1 _4386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4126__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2720_ _2789_/C _2718_/X _2706_/Y _2719_/Y vssd1 vssd1 vccd1 vccd1 _2720_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3965__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2651_ _4700_/Q vssd1 vssd1 vccd1 vccd1 _2651_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2582_ _4632_/Q vssd1 vssd1 vccd1 vccd1 _2722_/A sky130_fd_sc_hd__inv_2
X_4321_ _4080_/X _4421_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4321_/X sky130_fd_sc_hd__mux2_1
X_4252_ _4251_/X _4374_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4252_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3203_ _3234_/B _3198_/X _3152_/B vssd1 vssd1 vccd1 vccd1 _3204_/B sky130_fd_sc_hd__a21bo_1
X_4183_ _4183_/A vssd1 vssd1 vccd1 vccd1 _4183_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3134_ _3134_/A _3134_/B vssd1 vssd1 vccd1 vccd1 _3144_/A sky130_fd_sc_hd__or2_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3065_ _4545_/Q vssd1 vssd1 vccd1 vccd1 _3178_/A sky130_fd_sc_hd__inv_2
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3967_ _4767_/Q vssd1 vssd1 vccd1 vccd1 _3967_/Y sky130_fd_sc_hd__inv_2
X_2918_ _2918_/A vssd1 vssd1 vccd1 vccd1 _2918_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3898_ _4247_/X _4474_/Q _3900_/S vssd1 vssd1 vccd1 vccd1 _3899_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3594__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_30_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4558_/CLK sky130_fd_sc_hd__clkbuf_16
X_2849_ input5/X _2967_/A vssd1 vssd1 vccd1 vccd1 _2849_/X sky130_fd_sc_hd__or2_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4519_ _4589_/CLK _4519_/D vssd1 vssd1 vccd1 vccd1 _4519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4393__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4642_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4384__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2839__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3821_ _4510_/Q _3816_/X _4381_/X _3303_/A vssd1 vssd1 vccd1 vccd1 _4510_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4290__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4621_/CLK sky130_fd_sc_hd__clkbuf_16
X_3752_ _4561_/Q _3750_/X _2520_/A _3751_/X vssd1 vssd1 vccd1 vccd1 _4561_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3683_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3683_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2703_ _2703_/A _2703_/B vssd1 vssd1 vccd1 vccd1 _2704_/B sky130_fd_sc_hd__or2_1
X_2634_ _4646_/Q _4157_/A _4645_/Q _4156_/A vssd1 vssd1 vccd1 vccd1 _2636_/C sky130_fd_sc_hd__a22o_1
X_2565_ _4634_/Q _4145_/A _4635_/Q _2467_/A vssd1 vssd1 vccd1 vccd1 _2612_/B sky130_fd_sc_hd__o22a_1
X_4304_ _4303_/X _4429_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4304_/X sky130_fd_sc_hd__mux2_1
X_2496_ _2490_/X _2491_/X _2495_/X vssd1 vssd1 vccd1 vccd1 _2496_/X sky130_fd_sc_hd__a21bo_1
XFILLER_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4375__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4235_ _4234_/X _4370_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4235_/X sky130_fd_sc_hd__mux2_1
X_4166_ _4155_/A _4155_/B _4156_/B vssd1 vssd1 vccd1 vccd1 _4166_/X sky130_fd_sc_hd__a21bo_1
XFILLER_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3117_ _3117_/A _3117_/B vssd1 vssd1 vccd1 vccd1 _3118_/B sky130_fd_sc_hd__or2_1
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4097_ _4428_/X _4103_/B vssd1 vssd1 vccd1 vccd1 _4098_/A sky130_fd_sc_hd__and2_1
X_3048_ _4562_/Q vssd1 vssd1 vccd1 vccd1 _3051_/A sky130_fd_sc_hd__inv_2
XFILLER_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3246__A1 _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3797__A2 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3962__B _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2350_ _2255_/A _2255_/B _2318_/Y vssd1 vssd1 vccd1 vccd1 _2351_/B sky130_fd_sc_hd__a21o_1
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2281_ _2925_/A vssd1 vssd1 vccd1 vccd1 _3104_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4020_ _4020_/A _4039_/B _4020_/C vssd1 vssd1 vccd1 vccd1 _4020_/Y sky130_fd_sc_hd__nor3_2
Xclkbuf_leaf_1_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4744_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4285__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3237__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3804_ _4523_/Q _3802_/X _4394_/X _3800_/X vssd1 vssd1 vccd1 vccd1 _4523_/D sky130_fd_sc_hd__a22o_1
X_3735_ _3771_/A vssd1 vssd1 vccd1 vccd1 _3772_/A sky130_fd_sc_hd__inv_2
XANTENNA__4033__B _4033_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3666_ _4615_/Q _3600_/X _4237_/X _3602_/X vssd1 vssd1 vccd1 vccd1 _4615_/D sky130_fd_sc_hd__a22o_1
X_3597_ _3597_/A vssd1 vssd1 vccd1 vccd1 _4656_/D sky130_fd_sc_hd__clkbuf_1
X_2617_ _2616_/A _2568_/X _2611_/Y _2616_/X _2614_/X vssd1 vssd1 vccd1 vccd1 _2617_/X
+ sky130_fd_sc_hd__o221a_1
X_2548_ _2815_/A _2272_/B _2816_/A _2273_/A vssd1 vssd1 vccd1 vccd1 _2551_/B sky130_fd_sc_hd__o22a_1
XFILLER_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4218_ _4060_/X _4373_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4218_/X sky130_fd_sc_hd__mux2_1
X_2479_ input5/X _2487_/B input4/X _2355_/A vssd1 vssd1 vccd1 vccd1 _2489_/A sky130_fd_sc_hd__a22o_1
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4149_ _4149_/A _4149_/B vssd1 vssd1 vccd1 vccd1 _4150_/B sky130_fd_sc_hd__or2_1
XANTENNA__3228__A1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3779__A2 _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3951__A2 _3922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input46_A data_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3303__A _3303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2442__A2 _2377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3973__A _4094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3520_ _4354_/X _3556_/B _3594_/C vssd1 vssd1 vccd1 vccd1 _3536_/S sky130_fd_sc_hd__or3_4
X_3451_ _3451_/A vssd1 vssd1 vccd1 vccd1 _4722_/D sky130_fd_sc_hd__clkbuf_1
X_2402_ _4186_/X _2401_/B _3192_/A _2397_/B vssd1 vssd1 vccd1 vccd1 _2403_/D sky130_fd_sc_hd__a2bb2o_1
X_3382_ _3382_/A _3392_/B vssd1 vssd1 vccd1 vccd1 _4039_/C sky130_fd_sc_hd__or2_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2333_ _4598_/Q _2332_/Y _2273_/D vssd1 vssd1 vccd1 vccd1 _2334_/B sky130_fd_sc_hd__o21ai_1
XFILLER_97_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2264_ _4341_/X _2278_/A _2262_/X _2263_/Y vssd1 vssd1 vccd1 vccd1 _2306_/A sky130_fd_sc_hd__a22o_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4003_ _4208_/X _4007_/B vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__and2_1
XFILLER_92_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2969__B1 _2949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3630__A1 _4642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4767_ _4773_/CLK _4767_/D vssd1 vssd1 vccd1 vccd1 _4767_/Q sky130_fd_sc_hd__dfxtp_1
X_3718_ _3718_/A vssd1 vssd1 vccd1 vccd1 _3718_/X sky130_fd_sc_hd__clkbuf_2
X_4698_ _4750_/CLK _4698_/D vssd1 vssd1 vccd1 vccd1 _4698_/Q sky130_fd_sc_hd__dfxtp_1
X_3649_ _4629_/Q _3647_/X input3/X _3648_/X vssd1 vssd1 vccd1 vccd1 _4629_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3793__A _3814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3688__A1 _4602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2951_ _2951_/A _2951_/B vssd1 vssd1 vccd1 vccd1 _2951_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4621_ _4621_/CLK _4621_/D vssd1 vssd1 vccd1 vccd1 _4621_/Q sky130_fd_sc_hd__dfxtp_2
X_2882_ _2882_/A vssd1 vssd1 vccd1 vccd1 _2882_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4552_ _4556_/CLK _4552_/D vssd1 vssd1 vccd1 vccd1 _4552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4483_ _4706_/CLK _4483_/D vssd1 vssd1 vccd1 vccd1 _4483_/Q sky130_fd_sc_hd__dfxtp_1
X_3503_ _3503_/A vssd1 vssd1 vccd1 vccd1 _4697_/D sky130_fd_sc_hd__clkbuf_1
X_3434_ _4260_/X _4729_/Q _3442_/S vssd1 vssd1 vccd1 vccd1 _3435_/A sky130_fd_sc_hd__mux2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _3365_/A vssd1 vssd1 vccd1 vccd1 _3556_/B sky130_fd_sc_hd__buf_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _4343_/X vssd1 vssd1 vccd1 vccd1 _2317_/A sky130_fd_sc_hd__inv_2
X_3296_ _4770_/Q _3310_/B _3962_/A _3732_/C vssd1 vssd1 vccd1 vccd1 _4770_/D sky130_fd_sc_hd__o211a_1
X_2247_ _2247_/A _2247_/B vssd1 vssd1 vccd1 vccd1 _2248_/B sky130_fd_sc_hd__or2_1
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput79 _4524_/Q vssd1 vssd1 vccd1 vccd1 addr_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3788__A _3788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output77_A _4522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2333__A1 _4598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3150_ _3150_/A _3150_/B vssd1 vssd1 vccd1 vccd1 _3208_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3530__A0 _4284_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3081_ _3090_/A _3081_/B vssd1 vssd1 vccd1 vccd1 _3082_/B sky130_fd_sc_hd__or2_1
XFILLER_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4293__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3983_ _4201_/X _3995_/B vssd1 vssd1 vccd1 vccd1 _3984_/A sky130_fd_sc_hd__and2_1
X_2934_ _2292_/A _2928_/Y _4346_/X _2929_/Y _2933_/Y vssd1 vssd1 vccd1 vccd1 _2936_/C
+ sky130_fd_sc_hd__a221o_1
X_2865_ _4446_/Q vssd1 vssd1 vccd1 vccd1 _2995_/A sky130_fd_sc_hd__inv_2
X_4604_ _4695_/CLK _4604_/D vssd1 vssd1 vccd1 vccd1 _4604_/Q sky130_fd_sc_hd__dfxtp_2
X_4535_ _4571_/CLK _4535_/D vssd1 vssd1 vccd1 vccd1 _4535_/Q sky130_fd_sc_hd__dfxtp_1
X_2796_ _2737_/Y _2746_/X _2796_/C _2796_/D vssd1 vssd1 vccd1 vccd1 _2796_/X sky130_fd_sc_hd__and4bb_1
X_4466_ _4642_/CLK _4466_/D vssd1 vssd1 vccd1 vccd1 _4466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3417_ _3417_/A vssd1 vssd1 vccd1 vccd1 _4737_/D sky130_fd_sc_hd__clkbuf_1
X_4397_ _4637_/Q _4594_/Q _4559_/Q _4459_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4397_/X sky130_fd_sc_hd__mux4_1
XFILLER_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3348_ _3367_/A _3382_/A vssd1 vssd1 vccd1 vccd1 _4020_/C sky130_fd_sc_hd__or2_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3276_/A _3278_/X _3276_/B vssd1 vssd1 vccd1 vccd1 _3279_/X sky130_fd_sc_hd__o21ba_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2627__A2 _2536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3824__A1 _4507_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3824__B2 _3303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3760__B1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3815__A1 _4515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output115_A _4493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3815__B2 _3814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4240__A1 _3997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2650_ _2650_/A _2756_/A vssd1 vssd1 vccd1 vccd1 _2752_/B sky130_fd_sc_hd__or2_1
XFILLER_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2554__A1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3981__A _3981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2581_ _4633_/Q vssd1 vssd1 vccd1 vccd1 _2649_/A sky130_fd_sc_hd__inv_2
XFILLER_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4320_ _4319_/X _4422_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4320_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4251_ _4250_/X _4374_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4251_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4288__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3202_ _2412_/X _3197_/X _2409_/A _3201_/X vssd1 vssd1 vccd1 vccd1 _3210_/A sky130_fd_sc_hd__a22oi_1
X_4182_ _4145_/A _4145_/B _4146_/B vssd1 vssd1 vccd1 vccd1 _4182_/X sky130_fd_sc_hd__a21bo_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3133_ _3079_/A _3132_/X _3090_/D vssd1 vssd1 vccd1 vccd1 _3134_/B sky130_fd_sc_hd__a21bo_1
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3064_ _4548_/Q vssd1 vssd1 vccd1 vccd1 _3076_/A sky130_fd_sc_hd__inv_2
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3806__A1 _4521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2609__A2 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3806__B2 _3800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2490__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3966_ _3966_/A vssd1 vssd1 vccd1 vccd1 _3966_/X sky130_fd_sc_hd__clkbuf_1
X_2917_ _2266_/A _2911_/X _2912_/X _3033_/A vssd1 vssd1 vccd1 vccd1 _2937_/B sky130_fd_sc_hd__o211ai_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3897_ _3897_/A vssd1 vssd1 vccd1 vccd1 _4475_/D sky130_fd_sc_hd__clkbuf_1
X_2848_ _4448_/Q vssd1 vssd1 vccd1 vccd1 _2901_/A sky130_fd_sc_hd__inv_2
X_2779_ _2779_/A vssd1 vssd1 vccd1 vccd1 _2779_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3742__B1 _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4518_ _4518_/CLK _4518_/D vssd1 vssd1 vccd1 vccd1 _4518_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4198__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4449_ _4626_/CLK _4449_/D vssd1 vssd1 vccd1 vccd1 _4449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4393__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4289__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2210__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4384__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3041__A _3041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _4511_/Q _3816_/X _4382_/X _3814_/X vssd1 vssd1 vccd1 vccd1 _4511_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3751_ _3751_/A vssd1 vssd1 vccd1 vccd1 _3751_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2702_ _2702_/A _2702_/B vssd1 vssd1 vccd1 vccd1 _2703_/B sky130_fd_sc_hd__or2_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3682_ _3718_/A vssd1 vssd1 vccd1 vccd1 _3697_/A sky130_fd_sc_hd__buf_4
XFILLER_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2633_ _2668_/B _2537_/A _2668_/A _2816_/A vssd1 vssd1 vccd1 vccd1 _2638_/A sky130_fd_sc_hd__a22o_1
XANTENNA__3724__B1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2564_ _4638_/Q _4149_/A _4637_/Q _4148_/A vssd1 vssd1 vccd1 vccd1 _2616_/A sky130_fd_sc_hd__a22o_1
X_4303_ _4100_/X _4429_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4303_/X sky130_fd_sc_hd__mux2_1
X_2495_ _4114_/A _4578_/Q _2494_/X _4577_/Q vssd1 vssd1 vccd1 vccd1 _2495_/X sky130_fd_sc_hd__o22a_1
XFILLER_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4375__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4234_ _4052_/X _4370_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4234_/X sky130_fd_sc_hd__mux2_1
X_4165_ _4156_/A _4156_/B _4157_/B vssd1 vssd1 vccd1 vccd1 _4165_/X sky130_fd_sc_hd__a21bo_1
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3116_ _3116_/A _3119_/A vssd1 vssd1 vccd1 vccd1 _3117_/B sky130_fd_sc_hd__or2_1
X_4096_ _4096_/A vssd1 vssd1 vccd1 vccd1 _4096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3047_ _4563_/Q vssd1 vssd1 vccd1 vccd1 _3079_/A sky130_fd_sc_hd__inv_2
XFILLER_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_42_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3949_ _4442_/Q _3943_/X _2493_/A _3944_/X vssd1 vssd1 vccd1 vccd1 _4442_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3715__B1 _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2949__B _2949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2206__B1 _2204_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2205__A _2205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3706__B1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2280_ _4367_/X vssd1 vssd1 vccd1 vccd1 _2925_/A sky130_fd_sc_hd__inv_2
XFILLER_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2875__A _4456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2996__A1 _4447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3803_ _4524_/Q _3802_/X _4395_/X _3800_/X vssd1 vssd1 vccd1 vccd1 _4524_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3945__B1 _2505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3734_ _3750_/A vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3665_ _3665_/A vssd1 vssd1 vccd1 vccd1 _4616_/D sky130_fd_sc_hd__clkbuf_1
X_2616_ _2616_/A _2616_/B _2616_/C _2616_/D vssd1 vssd1 vccd1 vccd1 _2616_/X sky130_fd_sc_hd__or4_1
X_3596_ _4282_/X _4656_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3597_/A sky130_fd_sc_hd__mux2_1
X_2547_ _4157_/A _4603_/Q _4156_/A _4602_/Q vssd1 vssd1 vccd1 vccd1 _2549_/C sky130_fd_sc_hd__a22o_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2478_ input4/X _2355_/A _2471_/X _2477_/X vssd1 vssd1 vccd1 vccd1 _2478_/X sky130_fd_sc_hd__o211a_1
X_4217_ _4216_/X input35/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4217_/X sky130_fd_sc_hd__mux2_1
X_4148_ _4148_/A _4148_/B vssd1 vssd1 vccd1 vccd1 _4149_/B sky130_fd_sc_hd__or2_1
XFILLER_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4079_ _4421_/X _4081_/B vssd1 vssd1 vccd1 vccd1 _4080_/A sky130_fd_sc_hd__and2_1
XFILLER_43_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input39_A data_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_2_3_0_clk_A clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4416__A1 _4373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3927__B1 _2464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3450_ _4276_/X _4722_/Q _3458_/S vssd1 vssd1 vccd1 vccd1 _3451_/A sky130_fd_sc_hd__mux2_1
X_2401_ _4186_/X _2401_/B vssd1 vssd1 vccd1 vccd1 _2403_/C sky130_fd_sc_hd__and2_1
X_3381_ _3965_/A _3381_/B _4414_/X _3381_/D vssd1 vssd1 vccd1 vccd1 _3392_/B sky130_fd_sc_hd__or4_1
XFILLER_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2332_ _2332_/A _2332_/B vssd1 vssd1 vccd1 vccd1 _2332_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4296__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2263_ _2273_/A _2258_/B _2259_/B vssd1 vssd1 vccd1 vccd1 _2263_/Y sky130_fd_sc_hd__a21boi_1
X_4002_ _4038_/B _4006_/B vssd1 vssd1 vccd1 vccd1 _4002_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3918__B1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4766_ _4770_/CLK _4766_/D vssd1 vssd1 vccd1 vccd1 _4766_/Q sky130_fd_sc_hd__dfxtp_1
X_3717_ _3717_/A vssd1 vssd1 vccd1 vccd1 _3717_/X sky130_fd_sc_hd__clkbuf_2
X_4697_ _4742_/CLK _4697_/D vssd1 vssd1 vccd1 vccd1 _4697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3648_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3648_/X sky130_fd_sc_hd__buf_2
X_3579_ _4340_/X _4662_/Q _3606_/S vssd1 vssd1 vccd1 vccd1 _3580_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2950_ _2950_/A _2950_/B vssd1 vssd1 vccd1 vccd1 _2951_/B sky130_fd_sc_hd__or2_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ _2880_/A _2825_/X _2879_/Y _2824_/X _2880_/Y vssd1 vssd1 vccd1 vccd1 _2881_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4620_ _4621_/CLK _4620_/D vssd1 vssd1 vccd1 vccd1 _4620_/Q sky130_fd_sc_hd__dfxtp_1
X_4551_ _4583_/CLK _4551_/D vssd1 vssd1 vccd1 vccd1 _4551_/Q sky130_fd_sc_hd__dfxtp_1
X_4482_ _4701_/CLK _4482_/D vssd1 vssd1 vccd1 vccd1 _4482_/Q sky130_fd_sc_hd__dfxtp_1
X_3502_ _4260_/X _4697_/Q _3514_/S vssd1 vssd1 vccd1 vccd1 _3503_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3433_ _3728_/S vssd1 vssd1 vccd1 vccd1 _3442_/S sky130_fd_sc_hd__clkbuf_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4420__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3364_/A vssd1 vssd1 vccd1 vccd1 _3484_/A sky130_fd_sc_hd__buf_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3325_/B vssd1 vssd1 vccd1 vccd1 _3310_/B sky130_fd_sc_hd__inv_2
X_2315_ _2309_/A _2309_/B _2310_/B vssd1 vssd1 vccd1 vccd1 _2315_/X sky130_fd_sc_hd__a21bo_1
X_2246_ _2246_/A _2365_/A _2365_/B vssd1 vssd1 vccd1 vccd1 _2247_/B sky130_fd_sc_hd__or3_2
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4749_ _4750_/CLK _4749_/D vssd1 vssd1 vccd1 vccd1 _4749_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4411__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3833__S _3841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4402__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3080_ _3090_/B _3090_/D vssd1 vssd1 vccd1 vccd1 _3081_/B sky130_fd_sc_hd__or2_1
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _4033_/B _3994_/B vssd1 vssd1 vccd1 vccd1 _3982_/Y sky130_fd_sc_hd__nor2_1
X_2933_ _2933_/A vssd1 vssd1 vccd1 vccd1 _2933_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2864_ _4445_/Q vssd1 vssd1 vccd1 vccd1 _2994_/A sky130_fd_sc_hd__inv_2
X_4603_ _4695_/CLK _4603_/D vssd1 vssd1 vccd1 vccd1 _4603_/Q sky130_fd_sc_hd__dfxtp_2
X_2795_ _2789_/A _2720_/X _2786_/X _2798_/D _2794_/X vssd1 vssd1 vccd1 vccd1 _2799_/A
+ sky130_fd_sc_hd__o221a_1
X_4534_ _4571_/CLK _4534_/D vssd1 vssd1 vccd1 vccd1 _4534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4465_ _4565_/CLK _4465_/D vssd1 vssd1 vccd1 vccd1 _4465_/Q sky130_fd_sc_hd__dfxtp_1
X_3416_ _4288_/X _4737_/Q _3418_/S vssd1 vssd1 vccd1 vccd1 _3417_/A sky130_fd_sc_hd__mux2_1
X_4396_ _4636_/Q _4593_/Q _4558_/Q _4458_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4396_/X sky130_fd_sc_hd__mux4_2
X_3347_ _4014_/A _3366_/B vssd1 vssd1 vccd1 vccd1 _3382_/A sky130_fd_sc_hd__or2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3278_ _3275_/A _3277_/X _3275_/C vssd1 vssd1 vccd1 vccd1 _3278_/X sky130_fd_sc_hd__o21ba_1
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3824__A2 _3788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2229_ _2310_/A _2309_/A _2229_/C _2308_/A vssd1 vssd1 vccd1 vccd1 _2311_/B sky130_fd_sc_hd__or4_1
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3760__A1 _4555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2563__A2 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input21_A addr_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output108_A _4487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2580_ _2656_/A input3/X _2770_/A input2/X vssd1 vssd1 vccd1 vccd1 _2589_/B sky130_fd_sc_hd__a22o_1
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _4416_/X _4374_/X _4250_/S vssd1 vssd1 vccd1 vccd1 _4250_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3201_ _3076_/A _3076_/B _3196_/B vssd1 vssd1 vccd1 vccd1 _3201_/X sky130_fd_sc_hd__a21bo_1
X_4181_ _4181_/A vssd1 vssd1 vccd1 vccd1 _4181_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3132_ _3132_/A _3132_/B vssd1 vssd1 vccd1 vccd1 _3132_/X sky130_fd_sc_hd__or2_1
XANTENNA__3267__B1 _2543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3063_ _4549_/Q vssd1 vssd1 vccd1 vccd1 _3196_/A sky130_fd_sc_hd__inv_2
XANTENNA__3806__A2 _3802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2490__A1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3965_ _3965_/A _3965_/B _4773_/Q vssd1 vssd1 vccd1 vccd1 _3966_/A sky130_fd_sc_hd__or3_1
X_2916_ _2916_/A _2916_/B vssd1 vssd1 vccd1 vccd1 _3033_/A sky130_fd_sc_hd__or2_1
X_3896_ _4243_/X _4475_/Q _3896_/S vssd1 vssd1 vccd1 vccd1 _3897_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2847_ _4447_/Q vssd1 vssd1 vccd1 vccd1 _2896_/A sky130_fd_sc_hd__inv_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2778_ _2426_/A _2776_/B _2417_/A _2771_/X vssd1 vssd1 vccd1 vccd1 _2782_/C sky130_fd_sc_hd__a22o_1
X_4517_ _4518_/CLK _4517_/D vssd1 vssd1 vccd1 vccd1 _4517_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_clkbuf_leaf_1_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4448_ _4583_/CLK _4448_/D vssd1 vssd1 vccd1 vccd1 _4448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _4619_/Q _4576_/Q _4541_/Q _4441_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4379_/X sky130_fd_sc_hd__mux4_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3430__A0 _4256_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input69_A sb_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3497__B1 _4700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3249__B1 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4153__A _4153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3750_ _3750_/A vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2701_ _4210_/X _2698_/Y _2327_/X _2700_/Y vssd1 vssd1 vccd1 vccd1 _2709_/B sky130_fd_sc_hd__a22o_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3681_ _3717_/A vssd1 vssd1 vccd1 vccd1 _3718_/A sky130_fd_sc_hd__clkinv_4
X_2632_ _4643_/Q vssd1 vssd1 vccd1 vccd1 _2668_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__3724__B2 _3697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2527__A2 _4598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2563_ _2694_/A _2520_/A _2562_/X vssd1 vssd1 vccd1 vccd1 _2563_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4299__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4302_ _4301_/X _4430_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4302_/X sky130_fd_sc_hd__mux2_1
X_2494_ _2494_/A vssd1 vssd1 vccd1 vccd1 _2494_/X sky130_fd_sc_hd__clkbuf_2
X_4233_ _4232_/X _4005_/A _4354_/S vssd1 vssd1 vccd1 vccd1 _4233_/X sky130_fd_sc_hd__mux2_2
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4164_ _4157_/A _4157_/B _4158_/B vssd1 vssd1 vccd1 vccd1 _4164_/X sky130_fd_sc_hd__a21bo_1
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3115_ _3115_/A _3115_/B _3115_/C _3115_/D vssd1 vssd1 vccd1 vccd1 _3216_/D sky130_fd_sc_hd__or4_2
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4095_ _4369_/X _4103_/B vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__and2_1
XFILLER_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3046_ _4564_/Q vssd1 vssd1 vccd1 vccd1 _3090_/B sky130_fd_sc_hd__inv_2
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4047__B _4250_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3660__B1 _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3412__A0 _4284_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3948_ _4443_/Q _3943_/X _2492_/A _3944_/X vssd1 vssd1 vccd1 vccd1 _4443_/D sky130_fd_sc_hd__a22o_1
X_3879_ _4336_/X _4483_/Q _3885_/S vssd1 vssd1 vccd1 vccd1 _3880_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2311__A _2318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3841__S _3841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3651__B1 _2474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2206__B2 _3342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3052__A _4556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3642__B1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3802_ _3816_/A vssd1 vssd1 vccd1 vccd1 _3802_/X sky130_fd_sc_hd__buf_2
X_3733_ _3771_/A vssd1 vssd1 vccd1 vccd1 _3750_/A sky130_fd_sc_hd__buf_4
X_3664_ _4290_/X _4616_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3665_/A sky130_fd_sc_hd__mux2_1
X_2615_ _2702_/A input8/X _2614_/X vssd1 vssd1 vccd1 vccd1 _2616_/D sky130_fd_sc_hd__o21ai_1
X_3595_ _3958_/S vssd1 vssd1 vccd1 vccd1 _3780_/S sky130_fd_sc_hd__clkbuf_4
X_2546_ _2546_/A vssd1 vssd1 vccd1 vccd1 _4156_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2477_ input2/X _2418_/A _2474_/A _2413_/A _2476_/X vssd1 vssd1 vccd1 vccd1 _2477_/X
+ sky130_fd_sc_hd__o221a_1
X_4216_ _4016_/Y input35/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4216_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4147_ _4147_/A _4147_/B vssd1 vssd1 vccd1 vccd1 _4148_/B sky130_fd_sc_hd__or2_1
XFILLER_83_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3881__A0 _4338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4078_ _4078_/A vssd1 vssd1 vccd1 vccd1 _4078_/X sky130_fd_sc_hd__clkbuf_1
X_3029_ _3024_/A _2979_/Y _3011_/X _3041_/C _3028_/X vssd1 vssd1 vccd1 vccd1 _3029_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3624__B1 _2543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4416__A2 _4372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2400_ _2250_/A _2250_/B _2399_/Y vssd1 vssd1 vccd1 vccd1 _2401_/B sky130_fd_sc_hd__a21oi_1
X_3380_ _3380_/A vssd1 vssd1 vccd1 vccd1 _3381_/D sky130_fd_sc_hd__clkinv_2
X_2331_ _2953_/A vssd1 vssd1 vccd1 vccd1 _3134_/A sky130_fd_sc_hd__clkbuf_2
X_2262_ _2262_/A vssd1 vssd1 vccd1 vccd1 _2262_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_41_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4001_ _4001_/A vssd1 vssd1 vccd1 vccd1 _4038_/B sky130_fd_sc_hd__clkinv_2
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4765_ _4770_/CLK _4765_/D vssd1 vssd1 vccd1 vccd1 _4765_/Q sky130_fd_sc_hd__dfxtp_1
X_3716_ _4582_/Q _3710_/X _2507_/A _3711_/X vssd1 vssd1 vccd1 vccd1 _4582_/D sky130_fd_sc_hd__a22o_1
X_4696_ _4742_/CLK _4696_/D vssd1 vssd1 vccd1 vccd1 _4696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _3654_/A vssd1 vssd1 vccd1 vccd1 _3647_/X sky130_fd_sc_hd__buf_2
X_3578_ _4367_/S _3328_/A _3577_/Y _4663_/Q _3577_/A vssd1 vssd1 vccd1 vccd1 _4663_/D
+ sky130_fd_sc_hd__a32o_1
X_2529_ _2803_/A _2284_/A _2543_/A _2293_/A vssd1 vssd1 vccd1 vccd1 _2550_/A sky130_fd_sc_hd__a22o_1
XFILLER_88_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input51_A data_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4145__B _4145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ _2880_/A vssd1 vssd1 vccd1 vccd1 _2880_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _4583_/CLK _4550_/D vssd1 vssd1 vccd1 vccd1 _4550_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4481_ _4732_/CLK _4481_/D vssd1 vssd1 vccd1 vccd1 _4481_/Q sky130_fd_sc_hd__dfxtp_1
X_3501_ _3672_/S vssd1 vssd1 vccd1 vccd1 _3514_/S sky130_fd_sc_hd__clkbuf_4
X_3432_ _3484_/A _4353_/X _3588_/C vssd1 vssd1 vccd1 vccd1 _3728_/S sky130_fd_sc_hd__or3_4
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _3363_/A vssd1 vssd1 vccd1 vccd1 _4757_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4420__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2887__A1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _3121_/A _2314_/B vssd1 vssd1 vccd1 vccd1 _2433_/A sky130_fd_sc_hd__nor2_1
X_3294_ _4771_/Q _3291_/Y _2212_/X _3615_/B vssd1 vssd1 vccd1 vccd1 _4771_/D sky130_fd_sc_hd__o211a_1
X_2245_ _4576_/Q _4575_/Q _2244_/Y vssd1 vssd1 vccd1 vccd1 _2365_/B sky130_fd_sc_hd__o21ai_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4055__B _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4748_ _4750_/CLK _4748_/D vssd1 vssd1 vccd1 vccd1 _4748_/Q sky130_fd_sc_hd__dfxtp_1
X_4679_ _4733_/CLK _4679_/D vssd1 vssd1 vccd1 vccd1 _4679_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4411__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_51_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4732_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4402__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3325__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _3981_/A vssd1 vssd1 vccd1 vccd1 _4033_/B sky130_fd_sc_hd__clkinv_2
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2932_ _3110_/A _2932_/B vssd1 vssd1 vccd1 vccd1 _2933_/A sky130_fd_sc_hd__or2_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_42_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4771_/CLK sky130_fd_sc_hd__clkbuf_16
X_2863_ _2858_/X _2861_/X _2862_/X vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__a21bo_1
X_4602_ _4649_/CLK _4602_/D vssd1 vssd1 vccd1 vccd1 _4602_/Q sky130_fd_sc_hd__dfxtp_2
X_2794_ _2790_/Y _2791_/X _2690_/D _2689_/A _2793_/Y vssd1 vssd1 vccd1 vccd1 _2794_/X
+ sky130_fd_sc_hd__o32a_1
X_4533_ _4565_/CLK _4533_/D vssd1 vssd1 vccd1 vccd1 _4533_/Q sky130_fd_sc_hd__dfxtp_4
X_4464_ _4642_/CLK _4464_/D vssd1 vssd1 vccd1 vccd1 _4464_/Q sky130_fd_sc_hd__dfxtp_1
X_3415_ _3415_/A vssd1 vssd1 vccd1 vccd1 _4738_/D sky130_fd_sc_hd__clkbuf_1
X_4395_ _4635_/Q _4592_/Q _4557_/Q _4457_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4395_/X sky130_fd_sc_hd__mux4_2
XFILLER_97_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3346_ _3965_/A _3381_/B _4414_/X _3380_/A vssd1 vssd1 vccd1 vccd1 _3367_/A sky130_fd_sc_hd__or4_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3277_/A _3277_/B vssd1 vssd1 vccd1 vccd1 _3277_/X sky130_fd_sc_hd__and2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2228_ _4591_/Q vssd1 vssd1 vccd1 vccd1 _2308_/A sky130_fd_sc_hd__inv_2
XFILLER_26_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_33_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4719_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2548__B1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3844__S _3852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4396__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input14_A addr_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_24_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4638_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2539__B1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output82_A _4508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4387__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3200_ _2412_/X _3197_/X _2417_/X _3199_/X vssd1 vssd1 vccd1 vccd1 _3210_/B sky130_fd_sc_hd__o22ai_1
X_4180_ _4180_/A vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__clkbuf_1
X_3131_ _3130_/A _3132_/B _3137_/B vssd1 vssd1 vccd1 vccd1 _3131_/X sky130_fd_sc_hd__a21bo_1
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3267__A1 _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3062_ _4550_/Q vssd1 vssd1 vccd1 vccd1 _3198_/A sky130_fd_sc_hd__inv_2
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_15_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4518_/CLK sky130_fd_sc_hd__clkbuf_16
X_3964_ _4773_/Q vssd1 vssd1 vccd1 vccd1 _3964_/Y sky130_fd_sc_hd__inv_2
X_2915_ _4467_/Q _2907_/Y _2926_/B vssd1 vssd1 vccd1 vccd1 _2916_/B sky130_fd_sc_hd__o21ai_2
X_3895_ _3895_/A vssd1 vssd1 vccd1 vccd1 _4476_/D sky130_fd_sc_hd__clkbuf_1
X_2846_ _2482_/A _4455_/Q _2484_/A _4454_/Q _2845_/X vssd1 vssd1 vccd1 vccd1 _2851_/C
+ sky130_fd_sc_hd__a221o_1
X_2777_ _2409_/X _2773_/X _2783_/A _2776_/X vssd1 vssd1 vccd1 vccd1 _2782_/B sky130_fd_sc_hd__o211ai_1
XANTENNA__3664__S _3780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4516_ _4556_/CLK _4516_/D vssd1 vssd1 vccd1 vccd1 _4516_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4378__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4447_ _4583_/CLK _4447_/D vssd1 vssd1 vccd1 vccd1 _4447_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_input6_A addr_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4378_ _4618_/Q _4575_/Q _4540_/Q _4440_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4378_/X sky130_fd_sc_hd__mux4_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _4205_/X vssd1 vssd1 vccd1 vccd1 _3329_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3258__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3839__S _3841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3574__S _3606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4369__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3497__A1 _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3249__A1 _2500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2219__A _4599_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output120_A _4498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2700_ _2700_/A vssd1 vssd1 vccd1 vccd1 _2700_/Y sky130_fd_sc_hd__inv_2
X_3680_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3680_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2631_ _4642_/Q vssd1 vssd1 vccd1 vccd1 _2668_/B sky130_fd_sc_hd__inv_2
XANTENNA__3724__A2 _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2562_ _4641_/Q _2446_/A _2645_/C _2447_/A _2561_/X vssd1 vssd1 vccd1 vccd1 _2562_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4301_ _4102_/X _4430_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4301_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2493_ _2493_/A vssd1 vssd1 vccd1 vccd1 _2494_/A sky130_fd_sc_hd__inv_2
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4232_ _4008_/X _4005_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _4232_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4693_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4163_ _4158_/A _4158_/B _4159_/Y vssd1 vssd1 vccd1 vccd1 _4183_/A sky130_fd_sc_hd__a21oi_1
X_3114_ _3114_/A _3114_/B _3114_/C _3114_/D vssd1 vssd1 vccd1 vccd1 _3115_/D sky130_fd_sc_hd__or4_1
XFILLER_67_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4094_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4103_/B sky130_fd_sc_hd__buf_2
XFILLER_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3045_ _4565_/Q vssd1 vssd1 vccd1 vccd1 _3090_/A sky130_fd_sc_hd__inv_2
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3947_ _4444_/Q _3943_/X _2500_/A _3944_/X vssd1 vssd1 vccd1 vccd1 _4444_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2215__A2 _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3878_ _3878_/A vssd1 vssd1 vccd1 vccd1 _4484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2829_ _2456_/A _4459_/Q _2465_/A _4458_/Q vssd1 vssd1 vccd1 vccd1 _2874_/A sky130_fd_sc_hd__o22a_1
XANTENNA__2518__A3 _2510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3651__B2 _3648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3890__A1 _4478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_0_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3801_ _4525_/Q _3795_/X _4396_/X _3800_/X vssd1 vssd1 vccd1 vccd1 _4525_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3732_ _3965_/A _4771_/Q _3732_/C vssd1 vssd1 vccd1 vccd1 _3771_/A sky130_fd_sc_hd__or3_4
X_3663_ _4617_/Q _3600_/X _4241_/X _3602_/X vssd1 vssd1 vccd1 vccd1 _4617_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3508__A _3788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2614_ _4639_/Q _4150_/A _4638_/Q _2454_/A vssd1 vssd1 vccd1 vccd1 _2614_/X sky130_fd_sc_hd__o22a_1
X_3594_ _4354_/X _4353_/X _3594_/C vssd1 vssd1 vccd1 vccd1 _3958_/S sky130_fd_sc_hd__or3_4
X_2545_ _2545_/A vssd1 vssd1 vccd1 vccd1 _2546_/A sky130_fd_sc_hd__inv_2
X_2476_ _2473_/X _4583_/Q _2513_/A _4584_/Q vssd1 vssd1 vccd1 vccd1 _2476_/X sky130_fd_sc_hd__o22a_1
XFILLER_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4215_ _4214_/X input36/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4215_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4146_ _4146_/A _4146_/B vssd1 vssd1 vccd1 vccd1 _4147_/B sky130_fd_sc_hd__or2_1
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4077_ _4372_/X _4081_/B vssd1 vssd1 vccd1 vccd1 _4078_/A sky130_fd_sc_hd__and2_1
X_3028_ _3028_/A _3028_/B vssd1 vssd1 vccd1 vccd1 _3028_/X sky130_fd_sc_hd__or2_1
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3149__B1 _3119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3852__S _3852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ _4344_/X vssd1 vssd1 vccd1 vccd1 _2953_/A sky130_fd_sc_hd__inv_2
X_2261_ _4342_/X vssd1 vssd1 vccd1 vccd1 _2262_/A sky130_fd_sc_hd__inv_2
X_4000_ _4000_/A vssd1 vssd1 vccd1 vccd1 _4000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3863__A1 _4490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4764_ _4770_/CLK _4764_/D vssd1 vssd1 vccd1 vccd1 _4764_/Q sky130_fd_sc_hd__dfxtp_1
X_3715_ _4583_/Q _3710_/X _2472_/A _3711_/X vssd1 vssd1 vccd1 vccd1 _4583_/D sky130_fd_sc_hd__a22o_1
X_4695_ _4695_/CLK _4695_/D vssd1 vssd1 vccd1 vccd1 _4695_/Q sky130_fd_sc_hd__dfxtp_1
X_3646_ _4630_/Q _3640_/X input4/X _3641_/X vssd1 vssd1 vccd1 vccd1 _4630_/D sky130_fd_sc_hd__a22o_1
X_3577_ _3577_/A vssd1 vssd1 vccd1 vccd1 _3577_/Y sky130_fd_sc_hd__inv_2
X_2528_ _4152_/A _4598_/Q _2451_/Y _2525_/X _2527_/X vssd1 vssd1 vccd1 vccd1 _2528_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2459_ input8/X vssd1 vssd1 vccd1 vccd1 _2460_/A sky130_fd_sc_hd__inv_2
XFILLER_96_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4129_ _4129_/A _4129_/B vssd1 vssd1 vccd1 vccd1 _4130_/B sky130_fd_sc_hd__or2_1
XFILLER_56_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input44_A data_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4270__A1 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2227__A _4594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3058__A _4555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3500_ _4354_/X _3556_/B _3588_/C vssd1 vssd1 vccd1 vccd1 _3672_/S sky130_fd_sc_hd__or3_2
X_4480_ _4732_/CLK _4480_/D vssd1 vssd1 vccd1 vccd1 _4480_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2897__A _4661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3431_ _3431_/A vssd1 vssd1 vccd1 vccd1 _4730_/D sky130_fd_sc_hd__clkbuf_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _4229_/X _4757_/Q _3420_/S vssd1 vssd1 vccd1 vccd1 _3363_/A sky130_fd_sc_hd__mux2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2229_/C _2310_/X _2312_/Y vssd1 vssd1 vccd1 vccd1 _2314_/B sky130_fd_sc_hd__a21o_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3678_/A _3732_/C vssd1 vssd1 vccd1 vccd1 _3615_/B sky130_fd_sc_hd__or2_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2244_ _4665_/Q vssd1 vssd1 vccd1 vccd1 _2244_/Y sky130_fd_sc_hd__inv_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4747_ _4747_/CLK _4747_/D vssd1 vssd1 vccd1 vccd1 _4747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4678_ _4734_/CLK _4678_/D vssd1 vssd1 vccd1 vccd1 _4678_/Q sky130_fd_sc_hd__dfxtp_1
X_3629_ _4643_/Q _3626_/X _2816_/A _3627_/X vssd1 vssd1 vccd1 vccd1 _4643_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_40_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3763__B1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3818__A1 _4513_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3818__B2 _3814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3341__A _3341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _3980_/A vssd1 vssd1 vccd1 vccd1 _3980_/X sky130_fd_sc_hd__clkbuf_1
X_2931_ _4470_/Q _2922_/Y _2923_/X vssd1 vssd1 vccd1 vccd1 _2932_/B sky130_fd_sc_hd__o21ai_2
XFILLER_90_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_2862_ _4118_/A _4445_/Q _4117_/A _4444_/Q vssd1 vssd1 vccd1 vccd1 _2862_/X sky130_fd_sc_hd__o22a_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4601_ _4644_/CLK _4601_/D vssd1 vssd1 vccd1 vccd1 _4601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2793_ _2792_/X _2686_/A _2689_/B _2689_/D vssd1 vssd1 vccd1 vccd1 _2793_/Y sky130_fd_sc_hd__a31oi_2
X_4532_ _4644_/CLK _4532_/D vssd1 vssd1 vccd1 vccd1 _4532_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3754__B1 _2455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4463_ _4638_/CLK _4463_/D vssd1 vssd1 vccd1 vccd1 _4463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3414_ _4286_/X _4738_/Q _3418_/S vssd1 vssd1 vccd1 vccd1 _3415_/A sky130_fd_sc_hd__mux2_1
X_4394_ _4634_/Q _4591_/Q _4556_/Q _4456_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4394_/X sky130_fd_sc_hd__mux4_1
X_3345_ _4367_/S _4414_/X vssd1 vssd1 vccd1 vccd1 _3972_/A sky130_fd_sc_hd__nand2_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _3276_/A _3276_/B _3276_/C _3276_/D vssd1 vssd1 vccd1 vccd1 _3276_/X sky130_fd_sc_hd__or4_1
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _4594_/Q vssd1 vssd1 vccd1 vccd1 _2229_/C sky130_fd_sc_hd__inv_2
XFILLER_66_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4066__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2548__A1 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3745__B1 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4396__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2505__A _2505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2539__A1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4387__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output75_A _4520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4161__B1 _2536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3130_ _3130_/A _3132_/B vssd1 vssd1 vccd1 vccd1 _3137_/B sky130_fd_sc_hd__or2_1
X_3061_ _4551_/Q vssd1 vssd1 vccd1 vccd1 _3234_/B sky130_fd_sc_hd__inv_2
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4216__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3963_ _3963_/A vssd1 vssd1 vccd1 vccd1 _3963_/X sky130_fd_sc_hd__clkbuf_1
X_2914_ _2914_/A _2914_/B _2914_/C _2914_/D vssd1 vssd1 vccd1 vccd1 _2926_/B sky130_fd_sc_hd__or4_2
X_3894_ _4239_/X _4476_/Q _3896_/S vssd1 vssd1 vccd1 vccd1 _3895_/A sky130_fd_sc_hd__mux2_1
X_2845_ input7/X _2895_/A input6/X _2968_/A vssd1 vssd1 vccd1 vccd1 _2845_/X sky130_fd_sc_hd__a22o_1
X_4515_ _4556_/CLK _4515_/D vssd1 vssd1 vccd1 vccd1 _4515_/Q sky130_fd_sc_hd__dfxtp_2
X_2776_ _3204_/A _2776_/B vssd1 vssd1 vccd1 vccd1 _2776_/X sky130_fd_sc_hd__or2_1
X_4446_ _4623_/CLK _4446_/D vssd1 vssd1 vccd1 vccd1 _4446_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4378__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4377_ _4751_/Q _4702_/Q _4669_/Q _4612_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4377_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _3328_/A vssd1 vssd1 vccd1 vccd1 _4354_/S sky130_fd_sc_hd__buf_12
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3259_ _3237_/X _3244_/Y _3254_/X _3258_/X vssd1 vssd1 vccd1 vccd1 _3259_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__4077__A _4372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4207__A1 _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3855__S _3863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4369__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3497__A2 _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output113_A _4492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3041__D _3041_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2630_ _2667_/A _2545_/A _2667_/B _2815_/A vssd1 vssd1 vccd1 vccd1 _2636_/A sky130_fd_sc_hd__a22o_1
XANTENNA__3709__B1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2889__B _2889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2561_ _4640_/Q _2526_/A _2658_/A _2824_/A vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__o22a_1
X_2492_ _2492_/A vssd1 vssd1 vccd1 vccd1 _4114_/A sky130_fd_sc_hd__inv_2
X_4300_ _4299_/X _4431_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4300_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4231_ _4230_/X _4410_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4231_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4162_ _2532_/A _4159_/Y _4160_/X vssd1 vssd1 vccd1 vccd1 _4162_/Y sky130_fd_sc_hd__o21ai_1
X_3113_ _3104_/A _3104_/B _2301_/A _3110_/B vssd1 vssd1 vccd1 vccd1 _3114_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4093_ _4093_/A vssd1 vssd1 vccd1 vccd1 _4093_/X sky130_fd_sc_hd__clkbuf_1
X_3044_ _4566_/Q vssd1 vssd1 vccd1 vccd1 _3089_/B sky130_fd_sc_hd__inv_2
XFILLER_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3948__B1 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3946_ _4445_/Q _3943_/X _2498_/A _3944_/X vssd1 vssd1 vccd1 vccd1 _4445_/D sky130_fd_sc_hd__a22o_1
X_3877_ _4334_/X _4484_/Q _3885_/S vssd1 vssd1 vccd1 vccd1 _3878_/A sky130_fd_sc_hd__mux2_1
X_2828_ _2466_/A _4458_/Q _2467_/A _4457_/Q vssd1 vssd1 vccd1 vccd1 _2878_/B sky130_fd_sc_hd__a22o_1
X_2759_ _2762_/A _2762_/B _2390_/X _2758_/X vssd1 vssd1 vccd1 vccd1 _2765_/B sky130_fd_sc_hd__a22o_1
XFILLER_3_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4429_ _4743_/Q _4725_/Q _4692_/Q _4435_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4429_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3704__A _3718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3651__A2 _3647_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3939__B1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2850__B1 _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3800_ _3814_/A vssd1 vssd1 vccd1 vccd1 _3800_/X sky130_fd_sc_hd__buf_2
XFILLER_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3731_ _3731_/A vssd1 vssd1 vccd1 vccd1 _4572_/D sky130_fd_sc_hd__clkbuf_1
X_3662_ _4618_/Q _3633_/A input1/X _3634_/A vssd1 vssd1 vccd1 vccd1 _4618_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3593_ _3593_/A vssd1 vssd1 vccd1 vccd1 _4657_/D sky130_fd_sc_hd__clkbuf_1
X_2613_ _4634_/Q vssd1 vssd1 vccd1 vccd1 _2702_/A sky130_fd_sc_hd__inv_2
X_2544_ _2544_/A vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__clkbuf_2
X_2475_ _4130_/A vssd1 vssd1 vccd1 vccd1 _2513_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4214_ _4017_/Y input36/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4214_/X sky130_fd_sc_hd__mux2_1
X_4145_ _4145_/A _4145_/B vssd1 vssd1 vccd1 vccd1 _4146_/B sky130_fd_sc_hd__or2_1
XFILLER_95_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4076_ _4076_/A vssd1 vssd1 vccd1 vccd1 _4076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3027_ _3025_/C _3026_/Y _3020_/X vssd1 vssd1 vccd1 vccd1 _3028_/B sky130_fd_sc_hd__o21ai_1
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2841__B1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3929_ _3943_/A vssd1 vssd1 vccd1 vccd1 _3929_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3149__A1 _4555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4204__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4432__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2260_ _2272_/B _2259_/B _2259_/Y vssd1 vssd1 vccd1 vccd1 _2278_/A sky130_fd_sc_hd__a21oi_1
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4763_ _4771_/CLK _4763_/D vssd1 vssd1 vccd1 vccd1 _4763_/Q sky130_fd_sc_hd__dfxtp_1
X_3714_ _4584_/Q _3710_/X _2474_/A _3711_/X vssd1 vssd1 vccd1 vccd1 _4584_/D sky130_fd_sc_hd__a22o_1
X_4694_ _4752_/CLK _4694_/D vssd1 vssd1 vccd1 vccd1 _4694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4423__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3645_ _4631_/Q _3640_/X input5/X _3641_/X vssd1 vssd1 vccd1 vccd1 _4631_/D sky130_fd_sc_hd__a22o_1
X_3576_ _4354_/X _3576_/B _3581_/C vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__or3_1
X_2527_ _2446_/A _4598_/Q _4151_/A _4597_/Q vssd1 vssd1 vccd1 vccd1 _2527_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2458_ _4149_/A _4595_/Q _4148_/A _4594_/Q vssd1 vssd1 vccd1 vccd1 _2524_/A sky130_fd_sc_hd__a22o_1
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2389_ _4198_/X vssd1 vssd1 vccd1 vccd1 _2390_/A sky130_fd_sc_hd__inv_2
XFILLER_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4128_ input3/X vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__inv_2
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4059_ _4373_/X _4059_/B vssd1 vssd1 vccd1 vccd1 _4060_/A sky130_fd_sc_hd__and2_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2814__B1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3790__A1 _4533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3790__B2 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3863__S _3863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input37_A data_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3339__A _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4405__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3430_ _4256_/X _4730_/Q _3430_/S vssd1 vssd1 vccd1 vccd1 _3431_/A sky130_fd_sc_hd__mux2_1
X_3361_ _3361_/A vssd1 vssd1 vccd1 vccd1 _4758_/D sky130_fd_sc_hd__clkbuf_1
X_2312_ _2332_/B vssd1 vssd1 vccd1 vccd1 _2312_/Y sky130_fd_sc_hd__inv_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3292_ _4771_/Q vssd1 vssd1 vccd1 vccd1 _3678_/A sky130_fd_sc_hd__inv_2
X_2243_ _4577_/Q vssd1 vssd1 vccd1 vccd1 _2365_/A sky130_fd_sc_hd__inv_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4746_ _4746_/CLK _4746_/D vssd1 vssd1 vccd1 vccd1 _4746_/Q sky130_fd_sc_hd__dfxtp_1
X_4677_ _4735_/CLK _4677_/D vssd1 vssd1 vccd1 vccd1 _4677_/Q sky130_fd_sc_hd__dfxtp_1
X_3628_ _4644_/Q _3626_/X _2815_/A _3627_/X vssd1 vssd1 vccd1 vccd1 _4644_/D sky130_fd_sc_hd__a22o_1
X_3559_ _3559_/A vssd1 vssd1 vccd1 vccd1 _3560_/A sky130_fd_sc_hd__inv_2
XFILLER_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3818__A2 _3816_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ _2292_/X _2928_/Y _4346_/X _2929_/Y vssd1 vssd1 vccd1 vccd1 _2936_/B sky130_fd_sc_hd__o22ai_1
XFILLER_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ _2500_/A _2998_/A _2492_/A _2899_/A vssd1 vssd1 vccd1 vccd1 _2861_/X sky130_fd_sc_hd__o22a_1
X_4600_ _4600_/CLK _4600_/D vssd1 vssd1 vccd1 vccd1 _4600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2792_ _4347_/X _2792_/B vssd1 vssd1 vccd1 vccd1 _2792_/X sky130_fd_sc_hd__or2_1
X_4531_ _4531_/CLK _4531_/D vssd1 vssd1 vccd1 vccd1 _4531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4462_ _4565_/CLK _4462_/D vssd1 vssd1 vccd1 vccd1 _4462_/Q sky130_fd_sc_hd__dfxtp_1
X_3413_ _3413_/A vssd1 vssd1 vccd1 vccd1 _4739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4393_ _4633_/Q _4590_/Q _4555_/Q _4455_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4393_/X sky130_fd_sc_hd__mux4_1
X_3344_ _3349_/B vssd1 vssd1 vccd1 vccd1 _3974_/A sky130_fd_sc_hd__buf_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3275_ _3275_/A _3277_/A _3275_/C _3277_/B vssd1 vssd1 vccd1 vccd1 _3276_/D sky130_fd_sc_hd__or4b_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _4592_/Q vssd1 vssd1 vccd1 vccd1 _2309_/A sky130_fd_sc_hd__inv_2
XFILLER_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4729_ _4732_/CLK _4729_/D vssd1 vssd1 vccd1 vccd1 _4729_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4302__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4170__A1 _4153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3617__A _3633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4212__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4161__A1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3060_ _3060_/A _3148_/A vssd1 vssd1 vccd1 vccd1 _3078_/C sky130_fd_sc_hd__or2_1
XFILLER_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3672__A0 _4256_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3962_ _3962_/A _4338_/S _3962_/C vssd1 vssd1 vccd1 vccd1 _3963_/A sky130_fd_sc_hd__and3_1
X_2913_ _2913_/A _2913_/B vssd1 vssd1 vccd1 vccd1 _2914_/C sky130_fd_sc_hd__or2_1
X_3893_ _3893_/A vssd1 vssd1 vccd1 vccd1 _4477_/D sky130_fd_sc_hd__clkbuf_1
X_2844_ _4454_/Q vssd1 vssd1 vccd1 vccd1 _2968_/A sky130_fd_sc_hd__inv_2
XFILLER_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4514_ _4769_/CLK _4514_/D vssd1 vssd1 vccd1 vccd1 _4514_/Q sky130_fd_sc_hd__dfxtp_1
X_2775_ _2656_/A _2770_/X _2725_/B vssd1 vssd1 vccd1 vccd1 _2776_/B sky130_fd_sc_hd__a21bo_1
X_4445_ _4623_/CLK _4445_/D vssd1 vssd1 vccd1 vccd1 _4445_/Q sky130_fd_sc_hd__dfxtp_1
X_4376_ _4750_/Q _4701_/Q _4668_/Q _4610_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4376_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _3350_/A vssd1 vssd1 vccd1 vccd1 _3328_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3258_ input7/X _3060_/A _3240_/X _3257_/X vssd1 vssd1 vccd1 vccd1 _3258_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4077__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _4198_/X _3187_/A _3186_/Y _3188_/X vssd1 vssd1 vccd1 vccd1 _3193_/B sky130_fd_sc_hd__a211o_1
XFILLER_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2209_ _3299_/A vssd1 vssd1 vccd1 vccd1 _4338_/S sky130_fd_sc_hd__buf_12
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output106_A _4485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ _4641_/Q vssd1 vssd1 vccd1 vccd1 _2658_/A sky130_fd_sc_hd__inv_2
X_2491_ _2493_/A _2365_/A _3380_/A _2369_/Y vssd1 vssd1 vccd1 vccd1 _2491_/X sky130_fd_sc_hd__o22a_1
X_4230_ _4054_/X _4410_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4161_ _2532_/A _4159_/Y _2535_/A _2536_/X _4160_/X vssd1 vssd1 vccd1 vccd1 _4161_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3112_ _4351_/X _3219_/B _4346_/X _3107_/Y _3111_/Y vssd1 vssd1 vccd1 vccd1 _3114_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4092_ _4427_/X _4092_/B vssd1 vssd1 vccd1 vccd1 _4093_/A sky130_fd_sc_hd__and2_1
XFILLER_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3043_ _3043_/A _3042_/Y vssd1 vssd1 vccd1 vccd1 _3284_/A sky130_fd_sc_hd__or2b_1
XANTENNA__3645__B1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3945_ _4446_/Q _3943_/X _2505_/A _3944_/X vssd1 vssd1 vccd1 vccd1 _4446_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3876_ _3887_/A vssd1 vssd1 vccd1 vccd1 _3885_/S sky130_fd_sc_hd__buf_6
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2827_ _2460_/A _4456_/Q _2462_/A _4457_/Q vssd1 vssd1 vccd1 vccd1 _2874_/B sky130_fd_sc_hd__o22a_1
X_2758_ _2756_/A _2756_/B _2756_/Y vssd1 vssd1 vccd1 vccd1 _2758_/X sky130_fd_sc_hd__a21o_1
X_2689_ _2689_/A _2689_/B _2689_/C _2689_/D vssd1 vssd1 vccd1 vccd1 _2690_/D sky130_fd_sc_hd__or4_1
X_4428_ _4742_/Q _4724_/Q _4691_/Q _4651_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4428_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4359_ _4140_/X _4133_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4359_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3636__B1 _2452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3866__S _3874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input67_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4116__A1 _3381_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2850__A1 _2507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3730_ _4229_/X _4572_/Q _3730_/S vssd1 vssd1 vccd1 vccd1 _3731_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3661_ _4619_/Q _3633_/A _3380_/A _3634_/A vssd1 vssd1 vccd1 vccd1 _4619_/D sky130_fd_sc_hd__a22o_1
X_3592_ _4256_/X _4657_/Q _3952_/S vssd1 vssd1 vccd1 vccd1 _3593_/A sky130_fd_sc_hd__mux2_1
X_2612_ _2612_/A _2612_/B vssd1 vssd1 vccd1 vccd1 _2616_/C sky130_fd_sc_hd__nand2_1
X_2543_ _2543_/A vssd1 vssd1 vccd1 vccd1 _2544_/A sky130_fd_sc_hd__inv_2
X_2474_ _2474_/A vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__inv_2
X_4213_ _4212_/X input37/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4213_/X sky130_fd_sc_hd__mux2_2
X_4144_ _2472_/A _4121_/Y _4130_/B vssd1 vssd1 vccd1 vccd1 _4144_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4075_ _4420_/X _4081_/B vssd1 vssd1 vccd1 vccd1 _4076_/A sky130_fd_sc_hd__and2_1
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3026_ _3026_/A _3026_/B vssd1 vssd1 vccd1 vccd1 _3026_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2841__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3928_ _4457_/Q _3922_/X input9/X _3923_/X vssd1 vssd1 vccd1 vccd1 _4457_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4090__B _4092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3859_ _4318_/X _4492_/Q _3863_/S vssd1 vssd1 vccd1 vccd1 _3860_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4310__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3596__S _3780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4432__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4220__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4762_ _4771_/CLK _4762_/D vssd1 vssd1 vccd1 vccd1 _4762_/Q sky130_fd_sc_hd__dfxtp_1
X_3713_ _4585_/Q _3710_/X input2/X _3711_/X vssd1 vssd1 vccd1 vccd1 _4585_/D sky130_fd_sc_hd__a22o_1
X_4693_ _4693_/CLK _4693_/D vssd1 vssd1 vccd1 vccd1 _4693_/Q sky130_fd_sc_hd__dfxtp_1
X_3644_ _4632_/Q _3640_/X input6/X _3641_/X vssd1 vssd1 vccd1 vccd1 _4632_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4423__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3575_ _3575_/A vssd1 vssd1 vccd1 vccd1 _4664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2526_ _2526_/A vssd1 vssd1 vccd1 vccd1 _4151_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2457_ _2457_/A vssd1 vssd1 vccd1 vccd1 _4148_/A sky130_fd_sc_hd__clkbuf_1
X_2388_ _2248_/A _2248_/B _2249_/B vssd1 vssd1 vccd1 vccd1 _2393_/B sky130_fd_sc_hd__a21bo_1
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4127_ input4/X vssd1 vssd1 vccd1 vccd1 _4133_/A sky130_fd_sc_hd__inv_2
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4058_ _4058_/A vssd1 vssd1 vccd1 vccd1 _4058_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2814__A1 _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3009_ _3009_/A _3009_/B _3009_/C _3008_/X vssd1 vssd1 vccd1 vccd1 _3041_/A sky130_fd_sc_hd__or4b_2
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4305__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3790__A2 _3788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2805__A1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4215__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4405__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3355__A _3586_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output98_A _4512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3360_ _4225_/X _4758_/Q _3420_/S vssd1 vssd1 vccd1 vccd1 _3361_/A sky130_fd_sc_hd__mux2_1
X_2311_ _2318_/A _2311_/B vssd1 vssd1 vccd1 vccd1 _2332_/B sky130_fd_sc_hd__or2_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3732_/C vssd1 vssd1 vccd1 vccd1 _3291_/Y sky130_fd_sc_hd__inv_2
X_2242_ _4578_/Q vssd1 vssd1 vccd1 vccd1 _2246_/A sky130_fd_sc_hd__inv_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4751_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4745_ _4746_/CLK _4745_/D vssd1 vssd1 vccd1 vccd1 _4745_/Q sky130_fd_sc_hd__dfxtp_1
X_4676_ _4759_/CLK _4676_/D vssd1 vssd1 vccd1 vccd1 _4676_/Q sky130_fd_sc_hd__dfxtp_1
X_3627_ _3634_/A vssd1 vssd1 vccd1 vccd1 _3627_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3558_ _3559_/A vssd1 vssd1 vccd1 vccd1 _3558_/X sky130_fd_sc_hd__clkbuf_2
X_2509_ _2506_/X _4581_/Q _2508_/X _4582_/Q vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__o22a_1
X_3489_ _4706_/Q _3486_/X _4233_/X _3488_/X vssd1 vssd1 vccd1 vccd1 _4706_/D sky130_fd_sc_hd__a22o_1
XANTENNA__2648__D_N _4637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_36_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4734_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3874__S _3874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4399__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2723__B1 _2702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output136_A _2207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4738_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2860_ _4443_/Q vssd1 vssd1 vccd1 vccd1 _2899_/A sky130_fd_sc_hd__inv_2
XFILLER_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2791_ _2690_/A _2666_/X _2690_/C vssd1 vssd1 vccd1 vccd1 _2791_/X sky130_fd_sc_hd__o21ba_1
X_4530_ _4638_/CLK _4530_/D vssd1 vssd1 vccd1 vccd1 _4530_/Q sky130_fd_sc_hd__dfxtp_4
X_4461_ _4638_/CLK _4461_/D vssd1 vssd1 vccd1 vccd1 _4461_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3412_ _4284_/X _4739_/Q _3412_/S vssd1 vssd1 vccd1 vccd1 _3413_/A sky130_fd_sc_hd__mux2_1
X_4392_ _4632_/Q _4589_/Q _4554_/Q _4454_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4392_/X sky130_fd_sc_hd__mux4_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3965_/A _3366_/B vssd1 vssd1 vccd1 vccd1 _3349_/B sky130_fd_sc_hd__or2_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3274_ _2815_/A _3089_/B _2816_/A _3090_/A vssd1 vssd1 vccd1 vccd1 _3277_/B sky130_fd_sc_hd__o22a_1
XFILLER_58_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _4593_/Q vssd1 vssd1 vccd1 vccd1 _2310_/A sky130_fd_sc_hd__inv_2
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4649_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2989_ _2980_/A _2980_/B _2980_/Y vssd1 vssd1 vccd1 vccd1 _2992_/B sky130_fd_sc_hd__a21oi_1
X_4728_ _4732_/CLK _4728_/D vssd1 vssd1 vccd1 vccd1 _4728_/Q sky130_fd_sc_hd__dfxtp_1
X_4659_ _4734_/CLK _4659_/D vssd1 vssd1 vccd1 vccd1 _4659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3633__A _3633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _3961_/A vssd1 vssd1 vccd1 vccd1 _4435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2912_ _2266_/A _2911_/X _2262_/A _2909_/Y vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__o2bb2a_1
X_3892_ _4235_/X _4477_/Q _3896_/S vssd1 vssd1 vccd1 vccd1 _3893_/A sky130_fd_sc_hd__mux2_1
X_2843_ _4455_/Q vssd1 vssd1 vccd1 vccd1 _2895_/A sky130_fd_sc_hd__inv_2
X_2774_ _2412_/A _2769_/X _2409_/A _2773_/X vssd1 vssd1 vccd1 vccd1 _2783_/A sky130_fd_sc_hd__a22oi_1
X_4513_ _4625_/CLK _4513_/D vssd1 vssd1 vccd1 vccd1 _4513_/Q sky130_fd_sc_hd__dfxtp_2
X_4444_ _4623_/CLK _4444_/D vssd1 vssd1 vccd1 vccd1 _4444_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_7_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4589_/CLK sky130_fd_sc_hd__clkbuf_16
X_4375_ _4749_/Q _4699_/Q _4667_/Q _4609_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4375_/X sky130_fd_sc_hd__mux4_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _3904_/C vssd1 vssd1 vccd1 vccd1 _3350_/A sky130_fd_sc_hd__inv_2
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ input6/X _3148_/A _3244_/A _3256_/X _3242_/X vssd1 vssd1 vccd1 vccd1 _3257_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3188_ _2762_/A _3185_/B _2390_/X _3187_/Y vssd1 vssd1 vccd1 vccd1 _3188_/X sky130_fd_sc_hd__a22o_1
X_2208_ _3965_/B vssd1 vssd1 vccd1 vccd1 _3299_/A sky130_fd_sc_hd__inv_2
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3718__A _3718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4313__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input12_A addr_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2532__A _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4223__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3590__A0 _4264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2490_ _3380_/A _2369_/Y input1/X _2368_/Y vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__a211o_1
XANTENNA_output80_A _4525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4160_ _4160_/A _4160_/B vssd1 vssd1 vccd1 vccd1 _4160_/X sky130_fd_sc_hd__or2_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3111_ _3111_/A vssd1 vssd1 vccd1 vccd1 _3111_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4091_ _4091_/A vssd1 vssd1 vccd1 vccd1 _4091_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3042_ _3042_/A _3042_/B vssd1 vssd1 vccd1 vccd1 _3042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3944_ _3944_/A vssd1 vssd1 vccd1 vccd1 _3944_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3875_ _3875_/A vssd1 vssd1 vccd1 vccd1 _4485_/D sky130_fd_sc_hd__clkbuf_1
X_2826_ _2454_/A _4460_/Q _2457_/A _4459_/Q vssd1 vssd1 vccd1 vccd1 _2878_/A sky130_fd_sc_hd__a22o_1
XANTENNA__3538__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2757_ _4623_/Q _2756_/Y _2753_/B vssd1 vssd1 vccd1 vccd1 _2762_/B sky130_fd_sc_hd__o21ai_1
X_2688_ _2925_/A _2678_/B _2301_/A _2685_/B vssd1 vssd1 vccd1 vccd1 _2689_/D sky130_fd_sc_hd__a22o_1
X_4427_ _4747_/Q _4722_/Q _4689_/Q _4436_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4427_/X sky130_fd_sc_hd__mux4_1
XANTENNA_input4_A addr_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4358_ _4142_/X _2512_/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4358_/X sky130_fd_sc_hd__mux2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4088__B _4092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4022_/Y input40/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4289_/X sky130_fd_sc_hd__mux2_1
X_3309_ _3308_/Y _3306_/A _4767_/Q _3306_/Y vssd1 vssd1 vccd1 vccd1 _4767_/D sky130_fd_sc_hd__o22a_1
XFILLER_73_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3636__A1 _4638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4308__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3448__A _3484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4116__A2 _4013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4218__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3660_ _4620_/Q _3654_/X _2493_/A _3655_/X vssd1 vssd1 vccd1 vccd1 _4620_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3591_ _3591_/A vssd1 vssd1 vccd1 vccd1 _4658_/D sky130_fd_sc_hd__clkbuf_1
X_2611_ _2577_/X _2589_/Y _2606_/X _2610_/X vssd1 vssd1 vccd1 vccd1 _2611_/Y sky130_fd_sc_hd__a31oi_4
X_2542_ _2537_/A _2273_/B _2816_/A _2273_/A vssd1 vssd1 vccd1 vccd1 _2551_/A sky130_fd_sc_hd__a22o_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2473_ _4129_/A vssd1 vssd1 vccd1 vccd1 _2473_/X sky130_fd_sc_hd__clkbuf_2
X_4212_ _4018_/Y input37/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4212_/X sky130_fd_sc_hd__mux2_1
X_4143_ _2513_/X _4130_/B _4131_/B vssd1 vssd1 vccd1 vccd1 _4143_/X sky130_fd_sc_hd__a21bo_1
XFILLER_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4074_ _4074_/A vssd1 vssd1 vccd1 vccd1 _4074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3025_ _3026_/B _3025_/B _3025_/C _3028_/A vssd1 vssd1 vccd1 vccd1 _3041_/C sky130_fd_sc_hd__or4_2
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3927_ _4458_/Q _3922_/X _2464_/A _3923_/X vssd1 vssd1 vccd1 vccd1 _4458_/D sky130_fd_sc_hd__a22o_1
X_3858_ _3858_/A vssd1 vssd1 vccd1 vccd1 _4493_/D sky130_fd_sc_hd__clkbuf_1
X_3789_ _4534_/Q _3788_/X _4405_/X _3786_/X vssd1 vssd1 vccd1 vccd1 _4534_/D sky130_fd_sc_hd__a22o_1
X_2809_ _2535_/A _2806_/Y _2537_/A _2914_/B _2882_/A vssd1 vssd1 vccd1 vccd1 _2809_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3857__A1 _4493_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3877__S _3885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3906__A _3922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2810__A _4467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3641__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4273__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4761_ _4771_/CLK _4761_/D vssd1 vssd1 vccd1 vccd1 _4761_/Q sky130_fd_sc_hd__dfxtp_1
X_3712_ _4586_/Q _3710_/X input3/X _3711_/X vssd1 vssd1 vccd1 vccd1 _4586_/D sky130_fd_sc_hd__a22o_1
X_4692_ _4752_/CLK _4692_/D vssd1 vssd1 vccd1 vccd1 _4692_/Q sky130_fd_sc_hd__dfxtp_1
X_3643_ _4633_/Q _3640_/X input7/X _3641_/X vssd1 vssd1 vccd1 vccd1 _4633_/D sky130_fd_sc_hd__a22o_1
X_3574_ _4292_/X _4664_/Q _3606_/S vssd1 vssd1 vccd1 vccd1 _3575_/A sky130_fd_sc_hd__mux2_1
X_2525_ _2524_/A _2470_/X _2518_/Y _2524_/X _2522_/X vssd1 vssd1 vccd1 vccd1 _2525_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3839__A1 _4501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2456_ _2456_/A vssd1 vssd1 vccd1 vccd1 _2457_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2387_ _3185_/A vssd1 vssd1 vccd1 vccd1 _2762_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4126_ input5/X vssd1 vssd1 vccd1 vccd1 _4134_/A sky130_fd_sc_hd__inv_2
XFILLER_56_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4057_ _4415_/X _4059_/B vssd1 vssd1 vccd1 vccd1 _4058_/A sky130_fd_sc_hd__and2_1
XANTENNA__4264__A1 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3008_ _3008_/A _3008_/B vssd1 vssd1 vccd1 vccd1 _3008_/X sky130_fd_sc_hd__or2_1
XFILLER_71_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3775__B1 _2500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4321__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4255__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3766__B1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3230__A2 _4556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4231__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3290_/A _3325_/B vssd1 vssd1 vccd1 vccd1 _3732_/C sky130_fd_sc_hd__or2_1
X_2310_ _2310_/A _2310_/B vssd1 vssd1 vccd1 vccd1 _2310_/X sky130_fd_sc_hd__or2_1
X_2241_ _4579_/Q vssd1 vssd1 vccd1 vccd1 _2247_/A sky130_fd_sc_hd__inv_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3371__A _3484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4246__A1 _4375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4744_ _4744_/CLK _4744_/D vssd1 vssd1 vccd1 vccd1 _4744_/Q sky130_fd_sc_hd__dfxtp_1
X_4675_ _4759_/CLK _4675_/D vssd1 vssd1 vccd1 vccd1 _4675_/Q sky130_fd_sc_hd__dfxtp_1
X_3626_ _3633_/A vssd1 vssd1 vccd1 vccd1 _3626_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3557_ _3557_/A vssd1 vssd1 vccd1 vccd1 _3559_/A sky130_fd_sc_hd__buf_2
X_2508_ _4120_/A vssd1 vssd1 vccd1 vccd1 _2508_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_4_0_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3488_ _3488_/A vssd1 vssd1 vccd1 vccd1 _3488_/X sky130_fd_sc_hd__buf_2
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2439_ _2435_/Y _2436_/X _2306_/D _2305_/A _2438_/Y vssd1 vssd1 vccd1 vccd1 _2439_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _4434_/X _4109_/B vssd1 vssd1 vccd1 vccd1 _4110_/A sky130_fd_sc_hd__and2_1
XFILLER_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4316__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3748__B1 _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4399__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3890__S _3896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3920__B1 _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A data_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4228__A1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2535__A _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4226__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3739__B1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2790_ _2790_/A vssd1 vssd1 vccd1 vccd1 _2790_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3366__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4460_ _4638_/CLK _4460_/D vssd1 vssd1 vccd1 vccd1 _4460_/Q sky130_fd_sc_hd__dfxtp_1
X_4391_ _4631_/Q _4588_/Q _4553_/Q _4453_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4391_/X sky130_fd_sc_hd__mux4_1
X_3411_ _3411_/A vssd1 vssd1 vccd1 vccd1 _4740_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3911__B1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3342_ _3342_/A _3342_/B vssd1 vssd1 vccd1 vccd1 _3366_/B sky130_fd_sc_hd__or2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _2544_/A _4568_/Q _2546_/A _4567_/Q vssd1 vssd1 vccd1 vccd1 _3275_/C sky130_fd_sc_hd__a22o_1
XFILLER_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2224_/A _2336_/A _2328_/A vssd1 vssd1 vccd1 vccd1 _2332_/A sky130_fd_sc_hd__or3_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4219__A1 _4373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2988_ _2988_/A _2988_/B vssd1 vssd1 vccd1 vccd1 _2988_/X sky130_fd_sc_hd__and2_1
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4727_ _4752_/CLK _4727_/D vssd1 vssd1 vccd1 vccd1 _4727_/Q sky130_fd_sc_hd__dfxtp_1
X_4658_ _4732_/CLK _4658_/D vssd1 vssd1 vccd1 vccd1 _4658_/Q sky130_fd_sc_hd__dfxtp_1
X_3609_ _3609_/A vssd1 vssd1 vccd1 vccd1 _4652_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2705__A1 _4637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4589_ _4589_/CLK _4589_/D vssd1 vssd1 vccd1 vccd1 _4589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3885__S _3885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4161__A3 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3960_ _4270_/X _4435_/Q _3960_/S vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2911_ _2914_/B _2914_/D _2906_/B vssd1 vssd1 vccd1 vccd1 _2911_/X sky130_fd_sc_hd__a21bo_1
X_3891_ _3891_/A vssd1 vssd1 vccd1 vccd1 _4478_/D sky130_fd_sc_hd__clkbuf_1
X_2842_ input3/X _2902_/A input2/X _3014_/A vssd1 vssd1 vccd1 vccd1 _2851_/B sky130_fd_sc_hd__a22o_1
X_2773_ _2655_/A _2655_/B _2768_/B vssd1 vssd1 vccd1 vccd1 _2773_/X sky130_fd_sc_hd__a21bo_1
X_4512_ _4769_/CLK _4512_/D vssd1 vssd1 vccd1 vccd1 _4512_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4137__B1 _4145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4443_ _4621_/CLK _4443_/D vssd1 vssd1 vccd1 vccd1 _4443_/Q sky130_fd_sc_hd__dfxtp_1
X_4374_ _4748_/Q _4698_/Q _4666_/Q _4607_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4374_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _3965_/A _3325_/B vssd1 vssd1 vccd1 vccd1 _3904_/C sky130_fd_sc_hd__or2_1
X_3256_ input4/X _3152_/A _3244_/B _3255_/Y _3234_/X vssd1 vssd1 vccd1 vccd1 _3256_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _3297_/B _2207_/B _2206_/X vssd1 vssd1 vccd1 vccd1 _3965_/B sky130_fd_sc_hd__or3b_1
X_3187_ _3187_/A vssd1 vssd1 vccd1 vccd1 _3187_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3734__A _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3909__A _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2614__B1 _4638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output73_A _4518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3110_ _3110_/A _3110_/B vssd1 vssd1 vccd1 vccd1 _3111_/A sky130_fd_sc_hd__or2_1
X_4090_ _4426_/X _4092_/B vssd1 vssd1 vccd1 vccd1 _4091_/A sky130_fd_sc_hd__and2_1
XFILLER_95_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3041_ _3041_/A _3041_/B _3041_/C _3041_/D vssd1 vssd1 vccd1 vccd1 _3042_/B sky130_fd_sc_hd__or4_1
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3943_ _3943_/A vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3874_ _4332_/X _4485_/Q _3874_/S vssd1 vssd1 vccd1 vccd1 _3875_/A sky130_fd_sc_hd__mux2_1
X_2825_ _2447_/A _2891_/C _2520_/A _2941_/A _2824_/X vssd1 vssd1 vccd1 vccd1 _2825_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3538__B _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2756_ _2756_/A _2756_/B vssd1 vssd1 vccd1 vccd1 _2756_/Y sky130_fd_sc_hd__nor2_1
X_2687_ _2292_/X _2681_/Y _4346_/X _2682_/Y _2686_/Y vssd1 vssd1 vccd1 vccd1 _2689_/C
+ sky130_fd_sc_hd__a221o_1
X_4426_ _4746_/Q _4721_/Q _4688_/Q _4539_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4426_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _4181_/Y input9/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4357_/X sky130_fd_sc_hd__mux2_2
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4287_/X input41/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4288_/X sky130_fd_sc_hd__mux2_1
X_3308_ _3308_/A vssd1 vssd1 vccd1 vccd1 _3308_/Y sky130_fd_sc_hd__inv_2
X_3239_ input3/X _3234_/B input2/X _3198_/A vssd1 vssd1 vccd1 vccd1 _3244_/B sky130_fd_sc_hd__a22o_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4324__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3448__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2611__A3 _2606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output111_A _4490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2543__A _2543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4234__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3590_ _4264_/X _4658_/Q _3952_/S vssd1 vssd1 vccd1 vccd1 _3591_/A sky130_fd_sc_hd__mux2_1
X_2610_ _2649_/A input7/X _2583_/X _2609_/X vssd1 vssd1 vccd1 vccd1 _2610_/X sky130_fd_sc_hd__o22a_1
X_2541_ _2545_/A _2272_/A _2815_/A _2272_/B vssd1 vssd1 vccd1 vccd1 _2549_/A sky130_fd_sc_hd__a22o_1
X_2472_ _2472_/A vssd1 vssd1 vccd1 vccd1 _4129_/A sky130_fd_sc_hd__inv_2
X_4211_ _4178_/X _4147_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4211_/X sky130_fd_sc_hd__mux2_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4142_ _2512_/X _4131_/B _4132_/B vssd1 vssd1 vccd1 vccd1 _4142_/X sky130_fd_sc_hd__a21bo_1
XFILLER_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4073_ _4419_/X _4081_/B vssd1 vssd1 vccd1 vccd1 _4074_/A sky130_fd_sc_hd__and2_1
XFILLER_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3024_ _3024_/A _3024_/B _3024_/C _3024_/D vssd1 vssd1 vccd1 vccd1 _3028_/A sky130_fd_sc_hd__or4_1
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3926_ _4459_/Q _3922_/X _2455_/A _3923_/X vssd1 vssd1 vccd1 vccd1 _4459_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4426__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3857_ _4316_/X _4493_/Q _3863_/S vssd1 vssd1 vccd1 vccd1 _3858_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3788_ _3788_/A vssd1 vssd1 vccd1 vccd1 _3788_/X sky130_fd_sc_hd__clkbuf_4
X_2808_ _2533_/A _4470_/Q _2536_/A _4471_/Q vssd1 vssd1 vccd1 vccd1 _2882_/A sky130_fd_sc_hd__o22a_1
X_2739_ _2651_/Y _4619_/Q _2591_/Y _2590_/Y _2738_/X vssd1 vssd1 vccd1 vccd1 _2742_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4099__B _4103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4409_ _4649_/Q _4606_/Q _4571_/Q _4471_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4409_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4319__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4417__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3922__A _3922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4229__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4760_ _4760_/CLK _4760_/D vssd1 vssd1 vccd1 vccd1 _4760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3784__B2 _3303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4408__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3711_ _3718_/A vssd1 vssd1 vccd1 vccd1 _3711_/X sky130_fd_sc_hd__clkbuf_2
X_4691_ _4742_/CLK _4691_/D vssd1 vssd1 vccd1 vccd1 _4691_/Q sky130_fd_sc_hd__dfxtp_1
X_3642_ _4634_/Q _3640_/X input8/X _3641_/X vssd1 vssd1 vccd1 vccd1 _4634_/D sky130_fd_sc_hd__a22o_1
X_3573_ _3730_/S vssd1 vssd1 vccd1 vccd1 _3606_/S sky130_fd_sc_hd__clkbuf_4
X_2524_ _2524_/A _2524_/B _2524_/C _2524_/D vssd1 vssd1 vccd1 vccd1 _2524_/X sky130_fd_sc_hd__or4_1
X_2455_ _2455_/A vssd1 vssd1 vccd1 vccd1 _2456_/A sky130_fd_sc_hd__inv_2
X_2386_ _4188_/X vssd1 vssd1 vccd1 vccd1 _3185_/A sky130_fd_sc_hd__inv_2
XANTENNA__3832__A _3900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4125_ _2501_/X _4117_/B _4118_/B vssd1 vssd1 vccd1 vccd1 _4125_/X sky130_fd_sc_hd__a21bo_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4056_ _4056_/A vssd1 vssd1 vccd1 vccd1 _4056_/X sky130_fd_sc_hd__clkbuf_1
X_3007_ _3181_/A _2997_/B _3192_/A _3008_/B vssd1 vssd1 vccd1 vccd1 _3009_/C sky130_fd_sc_hd__a22o_1
XFILLER_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3909_ _3923_/A vssd1 vssd1 vccd1 vccd1 _3909_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3888__S _3896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2240_ _4580_/Q vssd1 vssd1 vccd1 vccd1 _2248_/A sky130_fd_sc_hd__inv_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3371__B _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4743_ _4752_/CLK _4743_/D vssd1 vssd1 vccd1 vccd1 _4743_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3509__B2 _3303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4674_ _4760_/CLK _4674_/D vssd1 vssd1 vccd1 vccd1 _4674_/Q sky130_fd_sc_hd__dfxtp_1
X_3625_ _4645_/Q _3617_/X _2545_/A _3620_/X vssd1 vssd1 vccd1 vccd1 _4645_/D sky130_fd_sc_hd__a22o_1
X_3556_ _4354_/X _3556_/B _3598_/C vssd1 vssd1 vccd1 vccd1 _3557_/A sky130_fd_sc_hd__or3_1
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2507_ _2507_/A vssd1 vssd1 vccd1 vccd1 _4120_/A sky130_fd_sc_hd__inv_2
X_3487_ _3487_/A vssd1 vssd1 vccd1 vccd1 _3488_/A sky130_fd_sc_hd__inv_2
X_2438_ _2437_/X _2302_/A _2305_/B _2305_/D vssd1 vssd1 vccd1 vccd1 _2438_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2369_ _4576_/Q vssd1 vssd1 vccd1 vccd1 _2369_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3693__B1 _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4108_ _4108_/A vssd1 vssd1 vccd1 vccd1 _4108_/X sky130_fd_sc_hd__clkbuf_1
X_4039_ _4039_/A _4039_/B _4039_/C vssd1 vssd1 vccd1 vccd1 _4039_/Y sky130_fd_sc_hd__nor3_1
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3737__A _3751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4332__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3684__B1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input35_A data_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3436__A0 _4264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2816__A _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4242__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3647__A _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4390_ _4630_/Q _4587_/Q _4552_/Q _4452_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4390_/X sky130_fd_sc_hd__mux4_1
X_3410_ _4282_/X _4740_/Q _3412_/S vssd1 vssd1 vccd1 vccd1 _3411_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3911__A1 _4470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3341_ _3341_/A vssd1 vssd1 vccd1 vccd1 _3342_/B sky130_fd_sc_hd__inv_2
XFILLER_97_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _2537_/A _3090_/B _2816_/A _3090_/A vssd1 vssd1 vccd1 vccd1 _3277_/A sky130_fd_sc_hd__a22o_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _4595_/Q vssd1 vssd1 vccd1 vccd1 _2328_/A sky130_fd_sc_hd__inv_2
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2478__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2987_ _2377_/Y _2986_/X _4194_/X _2985_/B _2988_/A vssd1 vssd1 vccd1 vccd1 _2988_/B
+ sky130_fd_sc_hd__o221ai_1
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4726_ _4744_/CLK _4726_/D vssd1 vssd1 vccd1 vccd1 _4726_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2461__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4657_ _4744_/CLK _4657_/D vssd1 vssd1 vccd1 vccd1 _4657_/Q sky130_fd_sc_hd__dfxtp_1
X_3608_ _4284_/X _4652_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3609_/A sky130_fd_sc_hd__mux2_1
X_4588_ _4634_/CLK _4588_/D vssd1 vssd1 vccd1 vccd1 _4588_/Q sky130_fd_sc_hd__dfxtp_2
X_3539_ _3554_/S vssd1 vssd1 vccd1 vccd1 _3548_/S sky130_fd_sc_hd__buf_2
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4327__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3657__B1 _2498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3930__A _3944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4237__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2910_ _4341_/X _2918_/A _2262_/X _2909_/Y vssd1 vssd1 vccd1 vccd1 _2937_/A sky130_fd_sc_hd__a22o_1
XFILLER_92_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3890_ _4231_/X _4478_/Q _3896_/S vssd1 vssd1 vccd1 vccd1 _3891_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2841_ input5/X _2967_/A input4/X _2971_/A vssd1 vssd1 vccd1 vccd1 _2851_/A sky130_fd_sc_hd__a22o_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2772_ _2412_/A _2769_/X _2417_/A _2771_/X vssd1 vssd1 vccd1 vccd1 _2783_/B sky130_fd_sc_hd__o22ai_1
X_4511_ _4623_/CLK _4511_/D vssd1 vssd1 vccd1 vccd1 _4511_/Q sky130_fd_sc_hd__dfxtp_1
X_4442_ _4621_/CLK _4442_/D vssd1 vssd1 vccd1 vccd1 _4442_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4137__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4373_ _4757_/Q _4707_/Q _4674_/Q _4572_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4373_/X sky130_fd_sc_hd__mux4_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _3287_/B _3320_/X _4764_/Q _3319_/A _2212_/X vssd1 vssd1 vccd1 vccd1 _4764_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3255_ _2512_/X _4550_/Q _2513_/A _4549_/Q _3235_/X vssd1 vssd1 vccd1 vccd1 _3255_/Y
+ sky130_fd_sc_hd__a221oi_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2202_/A _3287_/B _2204_/Y _3342_/A vssd1 vssd1 vccd1 vccd1 _2206_/X sky130_fd_sc_hd__a22o_1
X_3186_ _3186_/A vssd1 vssd1 vccd1 vccd1 _3186_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2871__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4709_ _4759_/CLK _4709_/D vssd1 vssd1 vccd1 vccd1 _4709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3750__A _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3639__B1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3896__S _3896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2614__A1 _4639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3811__B1 _4389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4367__A1 _2536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3040_ _2377_/Y _2986_/X _2988_/B _3039_/X vssd1 vssd1 vccd1 vccd1 _3041_/B sky130_fd_sc_hd__a211o_1
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _4447_/Q _3936_/X _2507_/A _3937_/X vssd1 vssd1 vccd1 vccd1 _4447_/D sky130_fd_sc_hd__a22o_1
X_3873_ _3873_/A vssd1 vssd1 vccd1 vccd1 _4486_/D sky130_fd_sc_hd__clkbuf_1
X_2824_ _2824_/A _2904_/A vssd1 vssd1 vccd1 vccd1 _2824_/X sky130_fd_sc_hd__or2_1
X_2755_ _3181_/A _2755_/B vssd1 vssd1 vccd1 vccd1 _2765_/A sky130_fd_sc_hd__nor2_1
X_2686_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2686_/Y sky130_fd_sc_hd__inv_2
X_4425_ _4745_/Q _4720_/Q _4687_/Q _4505_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4425_/X sky130_fd_sc_hd__mux4_1
X_4356_ _4137_/Y _4136_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4356_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2541__B1 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _4773_/Q _3306_/Y _4338_/S _4768_/Q _3306_/A vssd1 vssd1 vccd1 vccd1 _4768_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _4023_/Y input41/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4287_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3238_ input5/X _3242_/B input4/X _3152_/A vssd1 vssd1 vccd1 vccd1 _3244_/A sky130_fd_sc_hd__a22o_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _3169_/A vssd1 vssd1 vccd1 vccd1 _3169_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4340__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4380__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2824__A _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3655__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2540_ _2536_/X _4606_/Q _4153_/A _4599_/Q _2539_/X vssd1 vssd1 vccd1 vccd1 _2550_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4250__S _4250_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2471_ input3/X _2471_/B vssd1 vssd1 vccd1 vccd1 _2471_/X sky130_fd_sc_hd__or2_1
X_4210_ _4175_/Y _2520_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4210_/X sky130_fd_sc_hd__mux2_2
X_4141_ _4132_/A _4132_/B _4133_/B vssd1 vssd1 vccd1 vccd1 _4141_/X sky130_fd_sc_hd__a21bo_1
X_4072_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4081_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_95_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3023_ _2779_/X _2976_/X _2973_/X _2975_/X vssd1 vssd1 vccd1 vccd1 _3024_/C sky130_fd_sc_hd__o211ai_1
XANTENNA__4371__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3925_ _4460_/Q _3922_/X _2452_/A _3923_/X vssd1 vssd1 vccd1 vccd1 _4460_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4426__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3856_ _3856_/A vssd1 vssd1 vccd1 vccd1 _4494_/D sky130_fd_sc_hd__clkbuf_1
X_3787_ _4535_/Q _3508_/X _4406_/X _3786_/X vssd1 vssd1 vccd1 vccd1 _4535_/D sky130_fd_sc_hd__a22o_1
X_2807_ _4464_/Q vssd1 vssd1 vccd1 vccd1 _2914_/B sky130_fd_sc_hd__inv_2
X_2738_ _4700_/Q _4618_/Q vssd1 vssd1 vccd1 vccd1 _2738_/X sky130_fd_sc_hd__or2_1
X_4408_ _4648_/Q _4605_/Q _4570_/Q _4470_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4408_/X sky130_fd_sc_hd__mux4_2
X_2669_ _4645_/Q _2661_/Y _2679_/B vssd1 vssd1 vccd1 vccd1 _2670_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__3504__S _3514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4339_ _4019_/Y input38/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4339_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2644__A _4638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4335__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4417__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input65_A hit_dtlb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2808__B2 _4471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4245__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3710_ _3717_/A vssd1 vssd1 vccd1 vccd1 _3710_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3784__A2 _3508_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4690_ _4690_/CLK _4690_/D vssd1 vssd1 vccd1 vccd1 _4690_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4408__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3641_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3641_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3572_ _4354_/X _4353_/X _3572_/C vssd1 vssd1 vccd1 vccd1 _3730_/S sky130_fd_sc_hd__or3_2
XANTENNA__3385__A _3430_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2523_ input8/X _2308_/A _2522_/X vssd1 vssd1 vccd1 vccd1 _2524_/D sky130_fd_sc_hd__o21ai_1
X_2454_ _2454_/A vssd1 vssd1 vccd1 vccd1 _4149_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2385_ _2380_/Y _2382_/X _2441_/D _2441_/C vssd1 vssd1 vccd1 vccd1 _2385_/X sky130_fd_sc_hd__o211a_1
XFILLER_68_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4124_ _2499_/X _4118_/B _4119_/B vssd1 vssd1 vccd1 vccd1 _4124_/X sky130_fd_sc_hd__a21bo_1
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 addr_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_48_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4706_/CLK sky130_fd_sc_hd__clkbuf_16
X_4055_ _4368_/X _4059_/B vssd1 vssd1 vccd1 vccd1 _4056_/A sky130_fd_sc_hd__and2_1
X_3006_ _2995_/A _2995_/B _2995_/Y vssd1 vssd1 vccd1 vccd1 _3008_/B sky130_fd_sc_hd__a21o_1
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2464__A _2464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3224__A1 _2377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3908_ _3944_/A vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__buf_4
XFILLER_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3839_ _4300_/X _4501_/Q _3841_/S vssd1 vssd1 vccd1 vccd1 _3840_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_39_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4757_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2374__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4742_ _4742_/CLK _4742_/D vssd1 vssd1 vccd1 vccd1 _4742_/Q sky130_fd_sc_hd__dfxtp_1
X_4673_ _4756_/CLK _4673_/D vssd1 vssd1 vccd1 vccd1 _4673_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3509__A2 _3508_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3624_ _4646_/Q _3617_/X _2543_/A _3620_/X vssd1 vssd1 vccd1 vccd1 _4646_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3843__A _3900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3555_ _3555_/A vssd1 vssd1 vccd1 vccd1 _4674_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4182__A2 _4145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2506_ _4119_/A vssd1 vssd1 vccd1 vccd1 _2506_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3486_ _3487_/A vssd1 vssd1 vccd1 vccd1 _3486_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2437_ _4347_/X _2437_/B vssd1 vssd1 vccd1 vccd1 _2437_/X sky130_fd_sc_hd__or2_1
XFILLER_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2459__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2368_ _4575_/Q vssd1 vssd1 vccd1 vccd1 _2368_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3693__A1 _4599_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2299_ _3110_/A vssd1 vssd1 vccd1 vccd1 _2301_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4107_ _4433_/X _4109_/B vssd1 vssd1 vccd1 vccd1 _4108_/A sky130_fd_sc_hd__and2_1
X_4038_ _4039_/A _4038_/B _4039_/C vssd1 vssd1 vccd1 vccd1 _4038_/Y sky130_fd_sc_hd__nor3_2
XFILLER_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input28_A addr_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output96_A _4510_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3340_ _3365_/A vssd1 vssd1 vccd1 vccd1 _3576_/B sky130_fd_sc_hd__clkbuf_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3271_ _2545_/A _3089_/A _2815_/A _3089_/B vssd1 vssd1 vccd1 vccd1 _3275_/A sky130_fd_sc_hd__a22o_1
XFILLER_3_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _4596_/Q vssd1 vssd1 vccd1 vccd1 _2336_/A sky130_fd_sc_hd__inv_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2986_ _2897_/Y _2853_/Y _2983_/X vssd1 vssd1 vccd1 vccd1 _2986_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4725_ _4752_/CLK _4725_/D vssd1 vssd1 vccd1 vccd1 _4725_/Q sky130_fd_sc_hd__dfxtp_1
X_4656_ _4719_/CLK _4656_/D vssd1 vssd1 vccd1 vccd1 _4656_/Q sky130_fd_sc_hd__dfxtp_1
X_4587_ _4589_/CLK _4587_/D vssd1 vssd1 vccd1 vccd1 _4587_/Q sky130_fd_sc_hd__dfxtp_1
X_3607_ _3607_/A vssd1 vssd1 vccd1 vccd1 _4653_/D sky130_fd_sc_hd__clkbuf_1
Xinput70 stall_dcache vssd1 vssd1 vccd1 vccd1 _3297_/B sky130_fd_sc_hd__buf_2
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3538_ _4354_/X _3556_/B _3572_/C vssd1 vssd1 vccd1 vccd1 _3554_/S sky130_fd_sc_hd__or3_4
XFILLER_88_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_51_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3469_ _3469_/A vssd1 vssd1 vccd1 vccd1 _4714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2469__A2 _4594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3512__S _3514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2641__A2 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4343__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4394__A2 _4556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3422__S _3586_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2840_ _4453_/Q vssd1 vssd1 vccd1 vccd1 _2967_/A sky130_fd_sc_hd__inv_2
XANTENNA__4253__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4385__A2 _4547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2771_ _2770_/A _2770_/B _2770_/X vssd1 vssd1 vccd1 vccd1 _2771_/X sky130_fd_sc_hd__a21bo_1
X_4510_ _4769_/CLK _4510_/D vssd1 vssd1 vccd1 vccd1 _4510_/Q sky130_fd_sc_hd__dfxtp_4
X_4441_ _4695_/CLK _4441_/D vssd1 vssd1 vccd1 vccd1 _4441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _4736_/Q _4715_/Q _4682_/Q _4616_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4372_/X sky130_fd_sc_hd__mux4_2
XFILLER_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _3965_/A _3323_/B vssd1 vssd1 vccd1 vccd1 _4765_/D sky130_fd_sc_hd__nor2_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3254_ _3251_/X _3252_/X _3253_/X vssd1 vssd1 vccd1 vccd1 _3254_/X sky130_fd_sc_hd__a21bo_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2205_/A vssd1 vssd1 vccd1 vccd1 _3342_/A sky130_fd_sc_hd__clkinv_2
X_3185_ _3185_/A _3185_/B vssd1 vssd1 vccd1 vccd1 _3186_/A sky130_fd_sc_hd__or2_1
XFILLER_26_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3820__B2 _3814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2472__A _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2969_ _4455_/Q _2968_/Y _2949_/B vssd1 vssd1 vccd1 vccd1 _2970_/B sky130_fd_sc_hd__o21ai_1
X_4708_ _4759_/CLK _4708_/D vssd1 vssd1 vccd1 vccd1 _4708_/Q sky130_fd_sc_hd__dfxtp_1
X_4639_ _4639_/CLK _4639_/D vssd1 vssd1 vccd1 vccd1 _4639_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3103__A3 _4571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4338__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3811__A1 _4518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4248__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3941_ _4448_/Q _3936_/X _2472_/A _3937_/X vssd1 vssd1 vccd1 vccd1 _4448_/D sky130_fd_sc_hd__a22o_1
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3872_ _4330_/X _4486_/Q _3874_/S vssd1 vssd1 vccd1 vccd1 _3873_/A sky130_fd_sc_hd__mux2_1
X_2823_ _4463_/Q vssd1 vssd1 vccd1 vccd1 _2904_/A sky130_fd_sc_hd__inv_2
X_2754_ _4625_/Q _2753_/Y _2655_/B vssd1 vssd1 vccd1 vccd1 _2755_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2685_ _3110_/A _2685_/B vssd1 vssd1 vccd1 vccd1 _2686_/A sky130_fd_sc_hd__or2_1
XANTENNA__4012__A _4013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4424_ _4740_/Q _4719_/Q _4686_/Q _4656_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4424_/X sky130_fd_sc_hd__mux4_1
X_4355_ _4138_/X _4136_/B _4367_/S vssd1 vssd1 vccd1 vccd1 _4355_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2541__A1 _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _3306_/A vssd1 vssd1 vccd1 vccd1 _3306_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _4285_/X input42/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4286_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3237_ input4/X _3152_/A _3234_/X _3236_/X vssd1 vssd1 vccd1 vccd1 _3237_/X sky130_fd_sc_hd__o211a_1
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3168_ _3072_/Y _3164_/Y _3166_/X vssd1 vssd1 vccd1 vccd1 _3169_/A sky130_fd_sc_hd__o21ai_2
XFILLER_39_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3099_ _3102_/B vssd1 vssd1 vccd1 vccd1 _3099_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2377__A _2377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4285__A1 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4380__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input10_A addr_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2599__B2 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3936__A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2470_ _2519_/B _2524_/B _2519_/A vssd1 vssd1 vccd1 vccd1 _2470_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3720__B1 _2498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4140_ _4133_/A _4133_/B _4134_/B vssd1 vssd1 vccd1 vccd1 _4140_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__2523__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4071_ _4071_/A vssd1 vssd1 vccd1 vccd1 _4071_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3022_ _2426_/A _3020_/B _2417_/A _3015_/X vssd1 vssd1 vccd1 vccd1 _3025_/C sky130_fd_sc_hd__a22o_1
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4371__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3924_ _4461_/Q _3922_/X _2520_/A _3923_/X vssd1 vssd1 vccd1 vccd1 _4461_/D sky130_fd_sc_hd__a22o_1
X_3855_ _4314_/X _4494_/Q _3863_/S vssd1 vssd1 vccd1 vccd1 _3856_/A sky130_fd_sc_hd__mux2_1
X_2806_ _4471_/Q vssd1 vssd1 vccd1 vccd1 _2806_/Y sky130_fd_sc_hd__inv_2
X_3786_ _3814_/A vssd1 vssd1 vccd1 vccd1 _3786_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4200__A1 _3985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2737_ _4192_/X _2747_/B vssd1 vssd1 vccd1 vccd1 _2737_/Y sky130_fd_sc_hd__nor2_1
X_2668_ _2668_/A _2668_/B _2668_/C _2668_/D vssd1 vssd1 vccd1 vccd1 _2679_/B sky130_fd_sc_hd__or4_2
X_4407_ _4647_/Q _4604_/Q _4569_/Q _4469_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4407_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2599_ _2756_/A _2500_/A _2653_/A _2492_/A vssd1 vssd1 vccd1 vccd1 _2599_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3581__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _4337_/X _4371_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4338_/X sky130_fd_sc_hd__mux2_2
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4267__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4269_ _4034_/Y input51/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4269_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input2_A addr_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3778__B1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4351__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2450__B1 _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3950__B1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input58_A data_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3702__B1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4258__A1 _3981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2808__A2 _4470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3430__S _3430_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3769__B1 _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4261__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3640_ _3654_/A vssd1 vssd1 vccd1 vccd1 _3640_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3571_ _4367_/S _3328_/A _3570_/Y _4665_/Q _3570_/A vssd1 vssd1 vccd1 vccd1 _4665_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3941__B1 _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2522_ _4150_/A _4596_/Q _2454_/A _4595_/Q vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2453_ _2453_/A vssd1 vssd1 vccd1 vccd1 _2454_/A sky130_fd_sc_hd__clkbuf_2
X_2384_ _4187_/X _2384_/B vssd1 vssd1 vccd1 vccd1 _2441_/C sky130_fd_sc_hd__or2_1
XFILLER_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4123_ _2506_/X _4119_/B _4120_/B vssd1 vssd1 vccd1 vccd1 _4123_/X sky130_fd_sc_hd__a21bo_1
X_4054_ _4054_/A vssd1 vssd1 vccd1 vccd1 _4054_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4249__A1 _3989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 addr_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_6
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3005_ _4198_/X _3003_/A _3002_/Y _3004_/X vssd1 vssd1 vccd1 vccd1 _3009_/B sky130_fd_sc_hd__a211o_1
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3907_ _3943_/A vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__3576__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3838_ _3838_/A vssd1 vssd1 vccd1 vccd1 _4502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3769_ _4548_/Q _3764_/X _2472_/A _3765_/X vssd1 vssd1 vccd1 vccd1 _4548_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3932__B1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4346__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4256__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4741_ _4744_/CLK _4741_/D vssd1 vssd1 vccd1 vccd1 _4741_/Q sky130_fd_sc_hd__dfxtp_1
X_4672_ _4757_/CLK _4672_/D vssd1 vssd1 vccd1 vccd1 _4672_/Q sky130_fd_sc_hd__dfxtp_1
X_3623_ _4647_/Q _3617_/X _2803_/A _3620_/X vssd1 vssd1 vccd1 vccd1 _4647_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3914__B1 _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3554_ _4229_/X _4674_/Q _3554_/S vssd1 vssd1 vccd1 vccd1 _3555_/A sky130_fd_sc_hd__mux2_1
X_2505_ _2505_/A vssd1 vssd1 vccd1 vccd1 _4119_/A sky130_fd_sc_hd__inv_2
X_3485_ _3485_/A vssd1 vssd1 vccd1 vccd1 _3487_/A sky130_fd_sc_hd__clkbuf_2
X_2436_ _2306_/A _2268_/X _2306_/C vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__o21ba_1
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2367_ _4192_/X _2383_/B vssd1 vssd1 vccd1 vccd1 _2367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2298_ _4348_/X vssd1 vssd1 vccd1 vccd1 _3110_/A sky130_fd_sc_hd__inv_2
XFILLER_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4106_ _4106_/A vssd1 vssd1 vccd1 vccd1 _4106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4037_ _4039_/A _4037_/B _4039_/C vssd1 vssd1 vccd1 vccd1 _4037_/Y sky130_fd_sc_hd__nor3_1
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4397__A0 _4637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3944__A _3944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output89_A _4533_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3270_ _2536_/X _4571_/Q _2538_/A _4564_/Q _3269_/X vssd1 vssd1 vccd1 vccd1 _3276_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _4597_/Q vssd1 vssd1 vccd1 vccd1 _2224_/A sky130_fd_sc_hd__inv_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2985_ _4194_/X _2985_/B vssd1 vssd1 vccd1 vccd1 _2988_/A sky130_fd_sc_hd__nand2_1
X_4724_ _4742_/CLK _4724_/D vssd1 vssd1 vccd1 vccd1 _4724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4655_ _4756_/CLK _4655_/D vssd1 vssd1 vccd1 vccd1 _4655_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3854__A _3900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput60 data_in[5] vssd1 vssd1 vccd1 vccd1 _3997_/A sky130_fd_sc_hd__clkbuf_4
X_4586_ _4626_/CLK _4586_/D vssd1 vssd1 vccd1 vccd1 _4586_/Q sky130_fd_sc_hd__dfxtp_1
X_3606_ _4221_/X _4653_/Q _3606_/S vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__mux2_1
X_3537_ _3537_/A vssd1 vssd1 vccd1 vccd1 _4682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3468_ _4292_/X _4714_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3469_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2419_ _2418_/A _2418_/B _2418_/X vssd1 vssd1 vccd1 vccd1 _2419_/X sky130_fd_sc_hd__a21bo_1
X_3399_ _3399_/A vssd1 vssd1 vccd1 vccd1 _4746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4394__A3 _4456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3764__A _3771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input40_A data_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2617__B1 _2611_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4385__A3 _4447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2770_ _2770_/A _2770_/B vssd1 vssd1 vccd1 vccd1 _2770_/X sky130_fd_sc_hd__or2_1
X_4440_ _4618_/CLK _4440_/D vssd1 vssd1 vccd1 vccd1 _4440_/Q sky130_fd_sc_hd__dfxtp_1
X_4371_ _4758_/Q _4708_/Q _4675_/Q _4654_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4371_/X sky130_fd_sc_hd__mux4_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _3318_/Y _3320_/X _3321_/Y _2202_/A _3319_/A vssd1 vssd1 vccd1 vccd1 _3323_/B
+ sky130_fd_sc_hd__o32a_1
X_3253_ _2506_/X _4546_/Q _2508_/X _4547_/Q vssd1 vssd1 vccd1 vccd1 _3253_/X sky130_fd_sc_hd__o22a_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3184_ _4545_/Q _3182_/Y _3179_/B vssd1 vssd1 vccd1 vccd1 _3185_/B sky130_fd_sc_hd__o21ai_1
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2204_/A vssd1 vssd1 vccd1 vccd1 _2204_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__2856__B1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3820__A2 _3816_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2968_ _2968_/A _2968_/B vssd1 vssd1 vccd1 vccd1 _2968_/Y sky130_fd_sc_hd__nor2_1
X_4707_ _4757_/CLK _4707_/D vssd1 vssd1 vccd1 vccd1 _4707_/Q sky130_fd_sc_hd__dfxtp_1
X_2899_ _2899_/A _2980_/A _2980_/B vssd1 vssd1 vccd1 vccd1 _2998_/B sky130_fd_sc_hd__or3_2
X_4638_ _4638_/CLK _4638_/D vssd1 vssd1 vccd1 vccd1 _4638_/Q sky130_fd_sc_hd__dfxtp_2
X_4569_ _4571_/CLK _4569_/D vssd1 vssd1 vccd1 vccd1 _4569_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_1_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3272__B1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4354__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2838__B1 _2474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _4449_/Q _3936_/X _2474_/A _3937_/X vssd1 vssd1 vccd1 vccd1 _4449_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4264__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3871_ _3871_/A vssd1 vssd1 vccd1 vccd1 _4487_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_50_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2822_ _4461_/Q vssd1 vssd1 vccd1 vccd1 _2941_/A sky130_fd_sc_hd__inv_2
X_2753_ _2753_/A _2753_/B vssd1 vssd1 vccd1 vccd1 _2753_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3608__S _3780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2684_ _4648_/Q _2675_/Y _2676_/X vssd1 vssd1 vccd1 vccd1 _2685_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4012__B _4033_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4423_ _4739_/Q _4718_/Q _4685_/Q _4652_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4423_/X sky130_fd_sc_hd__mux4_1
X_4354_ _3971_/A _4771_/Q _4354_/S vssd1 vssd1 vccd1 vccd1 _4354_/X sky130_fd_sc_hd__mux2_8
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _3965_/A _4337_/S vssd1 vssd1 vccd1 vccd1 _3306_/A sky130_fd_sc_hd__or2_1
XFILLER_100_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _4024_/Y input42/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4285_/X sky130_fd_sc_hd__mux2_1
X_3236_ input2/X _3198_/A _2474_/A _3196_/A _3235_/X vssd1 vssd1 vccd1 vccd1 _3236_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3167_ _3072_/Y _4541_/Q _3164_/Y _3165_/Y _3166_/X vssd1 vssd1 vccd1 vccd1 _3170_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_82_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3098_ _3098_/A _3105_/A _3105_/B vssd1 vssd1 vccd1 vccd1 _3102_/B sky130_fd_sc_hd__or3_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2483__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_18_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4429__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4349__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3245__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2599__A2 _2500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3796__A1 _4529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3428__S _3430_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output71_A _4507_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4259__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4070_ _4418_/X _4070_/B vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__and2_1
XFILLER_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3021_ _2409_/X _3017_/X _3026_/A _3020_/X vssd1 vssd1 vccd1 vccd1 _3025_/B sky130_fd_sc_hd__o211ai_1
XFILLER_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3236__B1 _2474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3787__B2 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3923_ _3923_/A vssd1 vssd1 vccd1 vccd1 _3923_/X sky130_fd_sc_hd__clkbuf_2
X_3854_ _3900_/S vssd1 vssd1 vccd1 vccd1 _3863_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2805_ _2532_/A _2923_/A _2803_/X _2883_/A vssd1 vssd1 vccd1 vccd1 _2805_/X sky130_fd_sc_hd__o211a_1
X_3785_ _3785_/A vssd1 vssd1 vccd1 vccd1 _3814_/A sky130_fd_sc_hd__buf_2
X_2736_ _4621_/Q _2735_/Y _2756_/B vssd1 vssd1 vccd1 vccd1 _2747_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__4023__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2667_ _2667_/A _2667_/B vssd1 vssd1 vccd1 vccd1 _2668_/C sky130_fd_sc_hd__or2_1
X_4406_ _4646_/Q _4603_/Q _4568_/Q _4468_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4406_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2598_ _4621_/Q vssd1 vssd1 vccd1 vccd1 _2653_/A sky130_fd_sc_hd__inv_2
XANTENNA__3581__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4337_ _4063_/X _4371_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4337_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4268_ _4267_/X input52/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4268_/X sky130_fd_sc_hd__mux2_2
XFILLER_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3219_ _4351_/X _3219_/B vssd1 vssd1 vccd1 vccd1 _3219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4199_ _3990_/Y _3989_/A _4209_/S vssd1 vssd1 vccd1 vccd1 _4199_/X sky130_fd_sc_hd__mux2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3227__B1 _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3778__B2 _3751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3950__B2 _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3772__A _3772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3702__B2 _3697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4194__A1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3570_ _3570_/A vssd1 vssd1 vccd1 vccd1 _3570_/Y sky130_fd_sc_hd__inv_2
X_2521_ _2521_/A vssd1 vssd1 vccd1 vccd1 _4150_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3682__A _3718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2452_ _2452_/A vssd1 vssd1 vccd1 vccd1 _2453_/A sky130_fd_sc_hd__inv_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2383_ _4192_/X _2383_/B vssd1 vssd1 vccd1 vccd1 _2441_/D sky130_fd_sc_hd__nand2_1
XFILLER_96_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4122_ _2508_/X _4120_/B _4121_/Y vssd1 vssd1 vccd1 vccd1 _4122_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4053_ _4410_/X _4059_/B vssd1 vssd1 vccd1 vccd1 _4054_/A sky130_fd_sc_hd__and2_1
X_3004_ _3185_/A _3001_/B _2390_/A _3003_/Y vssd1 vssd1 vccd1 vccd1 _3004_/X sky130_fd_sc_hd__a22o_1
Xinput3 addr_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_6
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3906_ _3922_/A vssd1 vssd1 vccd1 vccd1 _3906_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3837_ _4298_/X _4502_/Q _3841_/S vssd1 vssd1 vccd1 vccd1 _3838_/A sky130_fd_sc_hd__mux2_1
X_3768_ _4549_/Q _3764_/X _2474_/A _3765_/X vssd1 vssd1 vccd1 vccd1 _4549_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2719_ _2709_/B _2708_/X _2709_/A vssd1 vssd1 vccd1 vccd1 _2719_/Y sky130_fd_sc_hd__a21oi_1
X_3699_ _4595_/Q _3696_/X _2452_/A _3697_/X vssd1 vssd1 vccd1 vccd1 _4595_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4362__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_2_0_clk_A clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input70_A stall_dcache vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3687__B1 _2543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4272__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4740_ _4740_/CLK _4740_/D vssd1 vssd1 vccd1 vccd1 _4740_/Q sky130_fd_sc_hd__dfxtp_1
X_4671_ _4755_/CLK _4671_/D vssd1 vssd1 vccd1 vccd1 _4671_/Q sky130_fd_sc_hd__dfxtp_1
X_3622_ _4648_/Q _3617_/X _2532_/A _3620_/X vssd1 vssd1 vccd1 vccd1 _4648_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3914__A1 _4467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3553_ _3553_/A vssd1 vssd1 vccd1 vccd1 _4675_/D sky130_fd_sc_hd__clkbuf_1
X_2504_ _2498_/A _2248_/A _2505_/A _2249_/A vssd1 vssd1 vccd1 vccd1 _2504_/X sky130_fd_sc_hd__o22a_1
X_3484_ _3484_/A _4353_/X _3598_/C vssd1 vssd1 vccd1 vccd1 _3485_/A sky130_fd_sc_hd__or3_1
X_2435_ _2435_/A vssd1 vssd1 vccd1 vccd1 _2435_/Y sky130_fd_sc_hd__inv_2
X_2366_ _4578_/Q _2365_/Y _2247_/B vssd1 vssd1 vccd1 vccd1 _2383_/B sky130_fd_sc_hd__o21ai_2
X_4105_ _4432_/X _4109_/B vssd1 vssd1 vccd1 vccd1 _4106_/A sky130_fd_sc_hd__and2_1
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2297_ _2292_/X _2295_/Y _4346_/X _2296_/Y vssd1 vssd1 vccd1 vccd1 _2305_/B sky130_fd_sc_hd__o22ai_2
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4036_ _4036_/A _4036_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4036_/Y sky130_fd_sc_hd__nor3_1
XFILLER_71_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3850__A0 _4310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4357__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4397__A1 _4594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4105__B _4109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3436__S _3442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _4598_/Q vssd1 vssd1 vccd1 vccd1 _2256_/A sky130_fd_sc_hd__inv_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4267__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2635__B2 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2984_ _2897_/Y _4441_/Q _2853_/Y _2852_/Y _2983_/X vssd1 vssd1 vccd1 vccd1 _2985_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4723_ _4744_/CLK _4723_/D vssd1 vssd1 vccd1 vccd1 _4723_/Q sky130_fd_sc_hd__dfxtp_1
X_4654_ _4759_/CLK _4654_/D vssd1 vssd1 vccd1 vccd1 _4654_/Q sky130_fd_sc_hd__dfxtp_1
X_4585_ _4626_/CLK _4585_/D vssd1 vssd1 vccd1 vccd1 _4585_/Q sky130_fd_sc_hd__dfxtp_1
Xinput50 data_in[25] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_2
Xinput61 data_in[6] vssd1 vssd1 vccd1 vccd1 _4001_/A sky130_fd_sc_hd__clkbuf_2
X_3605_ _3605_/A vssd1 vssd1 vccd1 vccd1 _4654_/D sky130_fd_sc_hd__clkbuf_1
X_3536_ _4290_/X _4682_/Q _3536_/S vssd1 vssd1 vccd1 vccd1 _3537_/A sky130_fd_sc_hd__mux2_1
X_3467_ _3482_/S vssd1 vssd1 vccd1 vccd1 _3476_/S sky130_fd_sc_hd__buf_2
X_2418_ _2418_/A _2418_/B vssd1 vssd1 vccd1 vccd1 _2418_/X sky130_fd_sc_hd__or2_1
X_3398_ _4278_/X _4746_/Q _3412_/S vssd1 vssd1 vccd1 vccd1 _3399_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2349_ _2349_/A vssd1 vssd1 vccd1 vccd1 _3150_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4019_ _4020_/A _4038_/B _4020_/C vssd1 vssd1 vccd1 vccd1 _4019_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__2626__B2 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A data_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _4753_/Q _4703_/Q _4670_/Q _4655_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4370_/X sky130_fd_sc_hd__mux4_1
X_3321_ _4764_/Q _3321_/B vssd1 vssd1 vccd1 vccd1 _3321_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3690__A _3697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _2498_/A _3178_/A _2505_/A _3179_/A vssd1 vssd1 vccd1 vccd1 _3252_/X sky130_fd_sc_hd__o22a_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2856__A1 _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3183_ _3182_/A _3182_/B _3182_/Y vssd1 vssd1 vccd1 vccd1 _3187_/A sky130_fd_sc_hd__a21oi_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _2203_/A vssd1 vssd1 vccd1 vccd1 _2207_/B sky130_fd_sc_hd__buf_2
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4026__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2967_ _2967_/A _2967_/B _2971_/B vssd1 vssd1 vccd1 vccd1 _2968_/B sky130_fd_sc_hd__or3_1
X_2898_ _4441_/Q _4440_/Q _2897_/Y vssd1 vssd1 vccd1 vccd1 _2980_/B sky130_fd_sc_hd__o21ai_1
X_4706_ _4706_/CLK _4706_/D vssd1 vssd1 vccd1 vccd1 _4706_/Q sky130_fd_sc_hd__dfxtp_1
X_4637_ _4637_/CLK _4637_/D vssd1 vssd1 vccd1 vccd1 _4637_/Q sky130_fd_sc_hd__dfxtp_2
X_4568_ _4571_/CLK _4568_/D vssd1 vssd1 vccd1 vccd1 _4568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3519_ _3519_/A vssd1 vssd1 vccd1 vccd1 _4690_/D sky130_fd_sc_hd__clkbuf_1
X_4499_ _4629_/CLK _4499_/D vssd1 vssd1 vccd1 vccd1 _4499_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4392__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3272__A1 _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clkbuf_opt_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _4531_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4383__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2838__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3870_ _4328_/X _4487_/Q _3874_/S vssd1 vssd1 vccd1 vccd1 _3871_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2821_ _4462_/Q vssd1 vssd1 vccd1 vccd1 _2891_/C sky130_fd_sc_hd__inv_2
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clk clkbuf_opt_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4623_/CLK sky130_fd_sc_hd__clkbuf_16
X_2752_ _2756_/B _2752_/B vssd1 vssd1 vccd1 vccd1 _2753_/B sky130_fd_sc_hd__or2_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4280__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2683_ _2292_/X _2681_/Y _4346_/X _2682_/Y vssd1 vssd1 vccd1 vccd1 _2689_/B sky130_fd_sc_hd__o22ai_2
X_4422_ _4738_/Q _4717_/Q _4684_/Q _4574_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4422_/X sky130_fd_sc_hd__mux4_2
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4353_ _4042_/Y _4770_/Q _4354_/S vssd1 vssd1 vccd1 vccd1 _4353_/X sky130_fd_sc_hd__mux2_8
X_3304_ _3965_/A _4769_/Q _3303_/X vssd1 vssd1 vccd1 vccd1 _4769_/D sky130_fd_sc_hd__a21o_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4284_ _4283_/X input43/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4284_/X sky130_fd_sc_hd__mux2_2
XFILLER_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3235_ _2473_/X _4548_/Q _2513_/A _4549_/Q vssd1 vssd1 vccd1 vccd1 _3235_/X sky130_fd_sc_hd__o22a_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4374__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3166_ _4663_/Q _4540_/Q vssd1 vssd1 vccd1 vccd1 _3166_/X sky130_fd_sc_hd__or2_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3097_ _4568_/Q vssd1 vssd1 vccd1 vccd1 _3105_/A sky130_fd_sc_hd__inv_2
XFILLER_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4429__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3999_ _4209_/X _4007_/B vssd1 vssd1 vccd1 vccd1 _4000_/A sky130_fd_sc_hd__and2_1
XFILLER_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4190__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4365__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3245__A1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3796__A2 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2849__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3020_ _3204_/A _3020_/B vssd1 vssd1 vccd1 vccd1 _3020_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_0_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4742_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4275__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3236__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3787__A2 _3508_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3922_ _3922_/A vssd1 vssd1 vccd1 vccd1 _3922_/X sky130_fd_sc_hd__clkbuf_2
X_3853_ _3853_/A vssd1 vssd1 vccd1 vccd1 _4495_/D sky130_fd_sc_hd__clkbuf_1
X_2804_ _2531_/A _4469_/Q _2544_/A _4468_/Q vssd1 vssd1 vccd1 vccd1 _2883_/A sky130_fd_sc_hd__o22a_1
X_3784_ _4536_/Q _3508_/X _4407_/X _3303_/X vssd1 vssd1 vccd1 vccd1 _4536_/D sky130_fd_sc_hd__a22o_1
X_2735_ _2735_/A _2735_/B vssd1 vssd1 vccd1 vccd1 _2735_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4023__B _4033_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2666_ _2266_/A _2665_/X _2262_/X _2663_/Y vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_99_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4405_ _4645_/Q _4602_/Q _4567_/Q _4467_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4405_/X sky130_fd_sc_hd__mux4_1
X_2597_ _4622_/Q vssd1 vssd1 vccd1 vccd1 _2756_/A sky130_fd_sc_hd__inv_2
X_4336_ _4335_/X _4412_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4336_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4267_ _4035_/Y input52/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4267_/X sky130_fd_sc_hd__mux2_1
X_4198_ _4125_/X _2501_/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4198_/X sky130_fd_sc_hd__mux2_1
X_3218_ _3115_/A _3087_/X _3115_/C vssd1 vssd1 vccd1 vccd1 _3218_/X sky130_fd_sc_hd__o21ba_1
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3149_ _4555_/Q _3148_/Y _3119_/A vssd1 vssd1 vccd1 vccd1 _3150_/B sky130_fd_sc_hd__o21ai_1
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3778__A2 _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2450__A2 _4598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3950__A2 _3922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3702__A2 _3696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output102_A _4516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2520_ _2520_/A vssd1 vssd1 vccd1 vccd1 _2521_/A sky130_fd_sc_hd__inv_2
X_2451_ _2520_/A _2336_/A _2450_/X vssd1 vssd1 vccd1 vccd1 _2451_/Y sky130_fd_sc_hd__o21ai_1
X_2382_ _4187_/X _2384_/B vssd1 vssd1 vccd1 vccd1 _2382_/X sky130_fd_sc_hd__and2_1
X_4121_ _4129_/B vssd1 vssd1 vccd1 vccd1 _4121_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4052_ _4052_/A vssd1 vssd1 vccd1 vccd1 _4052_/X sky130_fd_sc_hd__clkbuf_1
Xinput4 addr_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_8
X_3003_ _3003_/A vssd1 vssd1 vccd1 vccd1 _3003_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3905_ _3943_/A vssd1 vssd1 vccd1 vccd1 _3922_/A sky130_fd_sc_hd__buf_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3836_ _3836_/A vssd1 vssd1 vccd1 vccd1 _4503_/D sky130_fd_sc_hd__clkbuf_1
X_3767_ _4550_/Q _3764_/X input2/X _3765_/X vssd1 vssd1 vccd1 vccd1 _4550_/D sky130_fd_sc_hd__a22o_1
X_2718_ _2788_/A _2716_/Y _2717_/X vssd1 vssd1 vccd1 vccd1 _2718_/X sky130_fd_sc_hd__o21a_1
X_3698_ _4596_/Q _3696_/X _2520_/A _3697_/X vssd1 vssd1 vccd1 vccd1 _4596_/D sky130_fd_sc_hd__a22o_1
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2649_ _2649_/A _2722_/A vssd1 vssd1 vccd1 vccd1 _2657_/C sky130_fd_sc_hd__or2_1
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4319_ _4082_/X _4422_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4319_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input63_A data_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3687__A1 _4603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4670_ _4755_/CLK _4670_/D vssd1 vssd1 vccd1 vccd1 _4670_/Q sky130_fd_sc_hd__dfxtp_1
X_3621_ _4649_/Q _3617_/X _2535_/A _3620_/X vssd1 vssd1 vccd1 vccd1 _4649_/D sky130_fd_sc_hd__a22o_1
X_3552_ _4225_/X _4675_/Q _3554_/S vssd1 vssd1 vccd1 vccd1 _3553_/A sky130_fd_sc_hd__mux2_1
X_2503_ _2496_/X _2497_/X _2502_/X vssd1 vssd1 vccd1 vccd1 _2503_/X sky130_fd_sc_hd__a21bo_1
X_3483_ _3483_/A vssd1 vssd1 vccd1 vccd1 _4707_/D sky130_fd_sc_hd__clkbuf_1
X_2434_ _2434_/A _2434_/B _2434_/C vssd1 vssd1 vccd1 vccd1 _2443_/D sky130_fd_sc_hd__or3_1
X_2365_ _2365_/A _2365_/B vssd1 vssd1 vccd1 vccd1 _2365_/Y sky130_fd_sc_hd__nor2_1
X_4104_ _4104_/A vssd1 vssd1 vccd1 vccd1 _4104_/X sky130_fd_sc_hd__clkbuf_1
X_2296_ _2293_/A _2293_/B _2293_/Y vssd1 vssd1 vccd1 vccd1 _2296_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4029__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4035_ _4036_/A _4035_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4035_/Y sky130_fd_sc_hd__nor3_1
XFILLER_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3819_ _4512_/Q _3816_/X _4383_/X _3814_/X vssd1 vssd1 vccd1 vccd1 _4512_/D sky130_fd_sc_hd__a22o_1
XFILLER_79_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3841__A1 _4500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2580__B2 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2635__A2 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4283__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2983_ _4661_/Q _4440_/Q vssd1 vssd1 vccd1 vccd1 _2983_/X sky130_fd_sc_hd__or2_1
XFILLER_34_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4722_ _4747_/CLK _4722_/D vssd1 vssd1 vccd1 vccd1 _4722_/Q sky130_fd_sc_hd__dfxtp_1
Xinput40 data_in[16] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_2
X_4653_ _4759_/CLK _4653_/D vssd1 vssd1 vccd1 vccd1 _4653_/Q sky130_fd_sc_hd__dfxtp_1
Xinput51 data_in[26] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_2
X_4584_ _4626_/CLK _4584_/D vssd1 vssd1 vccd1 vccd1 _4584_/Q sky130_fd_sc_hd__dfxtp_2
X_3604_ _4225_/X _4654_/Q _3606_/S vssd1 vssd1 vccd1 vccd1 _3605_/A sky130_fd_sc_hd__mux2_1
Xinput62 data_in[7] vssd1 vssd1 vccd1 vccd1 _4005_/A sky130_fd_sc_hd__buf_2
X_3535_ _3535_/A vssd1 vssd1 vccd1 vccd1 _4683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3466_ _3484_/A _4353_/X _3572_/C vssd1 vssd1 vccd1 vccd1 _3482_/S sky130_fd_sc_hd__or3_4
XFILLER_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2417_ _2417_/A vssd1 vssd1 vccd1 vccd1 _2417_/X sky130_fd_sc_hd__clkbuf_2
X_3397_ _3397_/A vssd1 vssd1 vccd1 vccd1 _4747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2348_ _4356_/X vssd1 vssd1 vccd1 vccd1 _2349_/A sky130_fd_sc_hd__inv_2
XFILLER_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2279_ _3092_/A _2275_/B _2277_/Y _2278_/Y vssd1 vssd1 vccd1 vccd1 _2306_/C sky130_fd_sc_hd__a22o_1
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4018_ _4020_/A _4037_/B _4020_/C vssd1 vssd1 vccd1 vccd1 _4018_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__2626__A2 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3823__B2 _3303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4193__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3823__A1 _4508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3598__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2562__B2 _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A addr_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3578__B1 _4663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output94_A _4537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3320_ _3320_/A vssd1 vssd1 vccd1 vccd1 _3320_/X sky130_fd_sc_hd__clkbuf_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3248_/X _3249_/X _3250_/X vssd1 vssd1 vccd1 vccd1 _3251_/X sky130_fd_sc_hd__a21bo_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4278__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3182_ _3182_/A _3182_/B vssd1 vssd1 vccd1 vccd1 _3182_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2202_/A _3287_/B _2202_/C vssd1 vssd1 vccd1 vccd1 _2203_/A sky130_fd_sc_hd__and3_1
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2608__A2 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3805__A1 _4522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3805__B2 _3800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2966_ _3032_/C _2964_/X _2953_/Y _2965_/Y vssd1 vssd1 vccd1 vccd1 _2966_/X sky130_fd_sc_hd__o22a_1
X_2897_ _4661_/Q vssd1 vssd1 vccd1 vccd1 _2897_/Y sky130_fd_sc_hd__inv_2
X_4705_ _4755_/CLK _4705_/D vssd1 vssd1 vccd1 vccd1 _4705_/Q sky130_fd_sc_hd__dfxtp_1
X_4636_ _4637_/CLK _4636_/D vssd1 vssd1 vccd1 vccd1 _4636_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3336__A3 _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4567_ _4571_/CLK _4567_/D vssd1 vssd1 vccd1 vccd1 _4567_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3741__B1 _2543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4498_ _4701_/CLK _4498_/D vssd1 vssd1 vccd1 vccd1 _4498_/Q sky130_fd_sc_hd__dfxtp_2
X_3518_ _4274_/X _4690_/Q _3672_/S vssd1 vssd1 vccd1 vccd1 _3519_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4188__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3449_ _3464_/S vssd1 vssd1 vccd1 vccd1 _3458_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_76_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4392__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2480__B1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4221__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4288__A1 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4383__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output132_A _4480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4127__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2820_ _2445_/A _4463_/Q _2526_/A _4462_/Q vssd1 vssd1 vccd1 vccd1 _2880_/A sky130_fd_sc_hd__o22a_1
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2751_ _2751_/A vssd1 vssd1 vccd1 vccd1 _3181_/A sky130_fd_sc_hd__clkbuf_2
X_2682_ _2679_/A _2679_/B _2679_/Y vssd1 vssd1 vccd1 vccd1 _2682_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4421_ _4737_/Q _4716_/Q _4683_/Q _4472_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4421_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3723__B1 _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4352_ _4169_/A _4154_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4352_/X sky130_fd_sc_hd__mux2_1
X_3303_ _3303_/A vssd1 vssd1 vccd1 vccd1 _3303_/X sky130_fd_sc_hd__buf_2
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4283_ _4025_/Y input43/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4283_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4279__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3234_ input3/X _3234_/B vssd1 vssd1 vccd1 vccd1 _3234_/X sky130_fd_sc_hd__or2_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4374__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3165_ _4541_/Q vssd1 vssd1 vccd1 vccd1 _3165_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3096_ _4569_/Q vssd1 vssd1 vccd1 vccd1 _3098_/A sky130_fd_sc_hd__inv_2
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3998_ _4037_/B _4006_/B vssd1 vssd1 vccd1 vccd1 _3998_/Y sky130_fd_sc_hd__nor2_1
X_2949_ _2949_/A _2949_/B vssd1 vssd1 vccd1 vccd1 _2950_/B sky130_fd_sc_hd__or2_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4619_ _4695_/CLK _4619_/D vssd1 vssd1 vccd1 vccd1 _4619_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__2517__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3714__B1 _2474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3786__A _3814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3705__B1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3921_ _4462_/Q _3915_/X _2447_/A _3916_/X vssd1 vssd1 vccd1 vccd1 _4462_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3696__A _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4291__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3852_ _4312_/X _4495_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3853_/A sky130_fd_sc_hd__mux2_1
X_2803_ _2803_/A _2921_/A vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__or2_1
X_3783_ _4537_/Q _3508_/X _4408_/X _3303_/X vssd1 vssd1 vccd1 vccd1 _4537_/D sky130_fd_sc_hd__a22o_1
X_2734_ _2727_/X _2729_/X _2781_/B _2781_/D vssd1 vssd1 vccd1 vccd1 _2734_/Y sky130_fd_sc_hd__a31oi_1
X_2665_ _2668_/B _2668_/D _2660_/B vssd1 vssd1 vccd1 vccd1 _2665_/X sky130_fd_sc_hd__a21bo_1
X_2596_ _2592_/X _2594_/X _2595_/X vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__a21bo_1
X_4404_ _4644_/Q _4601_/Q _4566_/Q _4466_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4404_/X sky130_fd_sc_hd__mux4_1
X_4335_ _4065_/X _4412_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4335_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4266_ _4265_/X input53/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4266_/X sky130_fd_sc_hd__mux2_2
X_3217_ _3217_/A vssd1 vssd1 vccd1 vccd1 _3217_/Y sky130_fd_sc_hd__inv_2
X_4197_ _3994_/Y _3993_/A _4209_/S vssd1 vssd1 vccd1 vccd1 _4197_/X sky130_fd_sc_hd__mux2_1
X_3148_ _3148_/A _3148_/B vssd1 vssd1 vccd1 vccd1 _3148_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3079_ _3079_/A _3132_/A _3119_/B _3119_/A vssd1 vssd1 vccd1 vccd1 _3090_/D sky130_fd_sc_hd__or4_2
XANTENNA__3935__B1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4112__B1 _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3926__B1 _2455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2450_ _2445_/A _4598_/Q _2447_/A _2224_/A _2449_/X vssd1 vssd1 vccd1 vccd1 _2450_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2381_ _2365_/A _2365_/B _2365_/Y vssd1 vssd1 vccd1 vccd1 _2384_/B sky130_fd_sc_hd__a21oi_1
X_4120_ _4120_/A _4120_/B vssd1 vssd1 vccd1 vccd1 _4129_/B sky130_fd_sc_hd__or2_1
X_4051_ _4370_/X _4059_/B vssd1 vssd1 vccd1 vccd1 _4052_/A sky130_fd_sc_hd__and2_1
XANTENNA__4286__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 addr_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_6
X_3002_ _3002_/A vssd1 vssd1 vccd1 vccd1 _3002_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4406__A1 _4603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3904_ _4771_/Q _4770_/Q _3904_/C vssd1 vssd1 vccd1 vccd1 _3943_/A sky130_fd_sc_hd__or3_4
X_3835_ _4296_/X _4503_/Q _3841_/S vssd1 vssd1 vccd1 vccd1 _3836_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3917__B1 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3766_ _4551_/Q _3764_/X input3/X _3765_/X vssd1 vssd1 vccd1 vccd1 _4551_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2717_ _4363_/X _2705_/X _4211_/X _2710_/Y vssd1 vssd1 vccd1 vccd1 _2717_/X sky130_fd_sc_hd__o22a_1
X_3697_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__buf_2
XANTENNA__4050__A _4109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2648_ _2704_/A _2703_/A _2702_/A _4637_/Q vssd1 vssd1 vccd1 vccd1 _2691_/B sky130_fd_sc_hd__or4b_1
X_2579_ _2721_/A input5/X _2725_/A input4/X vssd1 vssd1 vccd1 vccd1 _2589_/A sky130_fd_sc_hd__a22o_1
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4318_ _4317_/X _4423_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4318_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4249_ _4248_/X _3989_/A _4354_/S vssd1 vssd1 vccd1 vccd1 _4249_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4196__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2592__C1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input56_A data_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3620_ _3634_/A vssd1 vssd1 vccd1 vccd1 _3620_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3551_ _3551_/A vssd1 vssd1 vccd1 vccd1 _4676_/D sky130_fd_sc_hd__clkbuf_1
X_2502_ _2499_/X _4580_/Q _2501_/X _4579_/Q vssd1 vssd1 vccd1 vccd1 _2502_/X sky130_fd_sc_hd__o22a_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3482_ _4229_/X _4707_/Q _3482_/S vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2433_ _2433_/A _2433_/B _2433_/C _2433_/D vssd1 vssd1 vccd1 vccd1 _2434_/B sky130_fd_sc_hd__or4_1
XFILLER_69_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2364_ _2358_/X _2407_/B _2407_/D vssd1 vssd1 vccd1 vccd1 _2364_/X sky130_fd_sc_hd__o21ba_1
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4103_ _4431_/X _4103_/B vssd1 vssd1 vccd1 vccd1 _4104_/A sky130_fd_sc_hd__and2_1
X_2295_ _2437_/B vssd1 vssd1 vccd1 vccd1 _2295_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4034_ _4036_/A _4034_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4034_/Y sky130_fd_sc_hd__nor3_1
XFILLER_92_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2405__A3 _2443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3818_ _4513_/Q _3816_/X _4384_/X _3814_/X vssd1 vssd1 vccd1 vccd1 _4513_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3749_ _4562_/Q _3743_/X _2447_/A _3744_/X vssd1 vssd1 vccd1 vccd1 _4562_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4410__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_16_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2580__A2 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4401__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2982_ _4192_/X _2991_/B vssd1 vssd1 vccd1 vccd1 _3039_/A sky130_fd_sc_hd__nor2_1
X_4721_ _4746_/CLK _4721_/D vssd1 vssd1 vccd1 vccd1 _4721_/Q sky130_fd_sc_hd__dfxtp_1
X_4652_ _4740_/CLK _4652_/D vssd1 vssd1 vccd1 vccd1 _4652_/Q sky130_fd_sc_hd__dfxtp_1
Xinput30 addr_in[7] vssd1 vssd1 vccd1 vccd1 _2507_/A sky130_fd_sc_hd__buf_6
X_3603_ _4655_/Q _3600_/X _4245_/X _3602_/X vssd1 vssd1 vccd1 vccd1 _4655_/D sky130_fd_sc_hd__a22o_1
Xinput63 data_in[8] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_4
Xinput41 data_in[17] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_4
X_4583_ _4583_/CLK _4583_/D vssd1 vssd1 vccd1 vccd1 _4583_/Q sky130_fd_sc_hd__dfxtp_2
Xinput52 data_in[27] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_2
X_3534_ _4288_/X _4683_/Q _3536_/S vssd1 vssd1 vccd1 vccd1 _3535_/A sky130_fd_sc_hd__mux2_1
X_3465_ _3465_/A vssd1 vssd1 vccd1 vccd1 _4715_/D sky130_fd_sc_hd__clkbuf_1
X_2416_ _4358_/X vssd1 vssd1 vccd1 vccd1 _2417_/A sky130_fd_sc_hd__inv_2
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3396_ _4276_/X _4747_/Q _3412_/S vssd1 vssd1 vccd1 vccd1 _3397_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2347_ _2433_/A _2325_/X _2434_/A _2345_/Y _2346_/Y vssd1 vssd1 vccd1 vccd1 _2347_/X
+ sky130_fd_sc_hd__o32a_1
X_2278_ _2278_/A vssd1 vssd1 vccd1 vccd1 _2278_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4017_ _4020_/A _4036_/B _4017_/C vssd1 vssd1 vccd1 vccd1 _4017_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__3823__A2 _3788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3598__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3119__A _3119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input19_A addr_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3578__A1 _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _2499_/X _4545_/Q _2501_/X _4544_/Q vssd1 vssd1 vccd1 vccd1 _3250_/X sky130_fd_sc_hd__o22a_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2587__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3181_ _3181_/A _3181_/B vssd1 vssd1 vccd1 vccd1 _3193_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _4766_/Q vssd1 vssd1 vccd1 vccd1 _2202_/C sky130_fd_sc_hd__inv_2
XFILLER_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4294__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3805__A2 _3802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2965_ _2956_/B _2955_/X _2956_/A vssd1 vssd1 vccd1 vccd1 _2965_/Y sky130_fd_sc_hd__a21oi_1
X_4704_ _4756_/CLK _4704_/D vssd1 vssd1 vccd1 vccd1 _4704_/Q sky130_fd_sc_hd__dfxtp_1
X_2896_ _2896_/A _2995_/A vssd1 vssd1 vccd1 vccd1 _2900_/C sky130_fd_sc_hd__or2_1
X_4635_ _4637_/CLK _4635_/D vssd1 vssd1 vccd1 vccd1 _4635_/Q sky130_fd_sc_hd__dfxtp_2
X_4566_ _4642_/CLK _4566_/D vssd1 vssd1 vccd1 vccd1 _4566_/Q sky130_fd_sc_hd__dfxtp_1
X_3517_ _3517_/A vssd1 vssd1 vccd1 vccd1 _4691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4497_ _4701_/CLK _4497_/D vssd1 vssd1 vccd1 vccd1 _4497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3448_ _3484_/A _4353_/X _3594_/C vssd1 vssd1 vccd1 vccd1 _3464_/S sky130_fd_sc_hd__or3_4
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _4753_/Q _3373_/X _4245_/X _3375_/X vssd1 vssd1 vccd1 vccd1 _4753_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2480__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2750_ _4186_/X vssd1 vssd1 vccd1 vccd1 _2751_/A sky130_fd_sc_hd__inv_2
X_2681_ _2792_/B vssd1 vssd1 vccd1 vccd1 _2681_/Y sky130_fd_sc_hd__inv_2
X_4420_ _4735_/Q _4714_/Q _4681_/Q _4664_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4420_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3982__A _4033_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4351_ _4183_/Y _4158_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4351_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4289__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3302_ _3785_/A vssd1 vssd1 vccd1 vccd1 _3303_/A sky130_fd_sc_hd__buf_2
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4282_ _4281_/X input45/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4282_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3260_/B _3263_/B _3260_/A vssd1 vssd1 vccd1 vccd1 _3233_/X sky130_fd_sc_hd__o21a_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3164_ _4540_/Q vssd1 vssd1 vccd1 vccd1 _3164_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3095_ _3092_/A _3092_/B _2277_/Y _3094_/Y vssd1 vssd1 vccd1 vccd1 _3115_/C sky130_fd_sc_hd__a22o_1
XANTENNA__3239__B1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3997_ _3997_/A vssd1 vssd1 vccd1 vccd1 _4037_/B sky130_fd_sc_hd__clkinv_2
X_2948_ _4210_/X _2945_/Y _2327_/A _2947_/Y vssd1 vssd1 vccd1 vccd1 _2956_/B sky130_fd_sc_hd__a22o_1
XFILLER_50_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4618_ _4618_/CLK _4618_/D vssd1 vssd1 vccd1 vccd1 _4618_/Q sky130_fd_sc_hd__dfxtp_1
X_2879_ _2878_/A _2830_/X _2873_/Y _2878_/X _2876_/X vssd1 vssd1 vccd1 vccd1 _2879_/Y
+ sky130_fd_sc_hd__o221ai_2
X_4549_ _4583_/CLK _4549_/D vssd1 vssd1 vccd1 vccd1 _4549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2658__D _2702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3116__B _3119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3650__B1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3920_ _4463_/Q _3915_/X _2824_/A _3916_/X vssd1 vssd1 vccd1 vccd1 _4463_/D sky130_fd_sc_hd__a22o_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3977__A _4032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3851_ _3851_/A vssd1 vssd1 vccd1 vccd1 _4496_/D sky130_fd_sc_hd__clkbuf_1
X_3782_ _4538_/Q _3508_/X _4409_/X _3303_/X vssd1 vssd1 vccd1 vccd1 _4538_/D sky130_fd_sc_hd__a22o_1
X_2802_ _4469_/Q vssd1 vssd1 vccd1 vccd1 _2921_/A sky130_fd_sc_hd__inv_2
XANTENNA__4197__A1 _3993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2733_ _2349_/A _2724_/B _2360_/X _2729_/B vssd1 vssd1 vccd1 vccd1 _2781_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2664_ _4341_/X _2672_/A _2262_/X _2663_/Y vssd1 vssd1 vccd1 vccd1 _2690_/A sky130_fd_sc_hd__a22o_1
X_2595_ _4621_/Q _4114_/A _4620_/Q _2494_/X vssd1 vssd1 vccd1 vccd1 _2595_/X sky130_fd_sc_hd__o22a_1
X_4403_ _4643_/Q _4600_/Q _4565_/Q _4465_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4403_/X sky130_fd_sc_hd__mux4_1
X_4334_ _4333_/X _4413_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4334_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4265_ _4036_/Y input53/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4265_/X sky130_fd_sc_hd__mux2_1
X_3216_ _3216_/A _3216_/B _3216_/C _3216_/D vssd1 vssd1 vccd1 vccd1 _3225_/D sky130_fd_sc_hd__or4_2
X_4196_ _4195_/X _3962_/C _4338_/S vssd1 vssd1 vccd1 vccd1 _4196_/X sky130_fd_sc_hd__mux2_8
X_3147_ _3242_/B _3151_/A _3152_/B vssd1 vssd1 vccd1 vccd1 _3148_/B sky130_fd_sc_hd__or3_1
XFILLER_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3078_ _3242_/B _3151_/A _3078_/C _3152_/B vssd1 vssd1 vccd1 vccd1 _3119_/A sky130_fd_sc_hd__or4_4
XANTENNA__3632__B1 _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3699__B1 _2452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4112__A1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3623__B1 _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2380_ _4194_/X _2378_/B _2379_/X vssd1 vssd1 vccd1 vccd1 _2380_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_96_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _4109_/B vssd1 vssd1 vccd1 vccd1 _4059_/B sky130_fd_sc_hd__buf_2
XFILLER_1_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 addr_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_6
X_3001_ _3185_/A _3001_/B vssd1 vssd1 vccd1 vccd1 _3002_/A sky130_fd_sc_hd__or2_1
XFILLER_76_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3500__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3903_ _3903_/A vssd1 vssd1 vccd1 vccd1 _4472_/D sky130_fd_sc_hd__clkbuf_1
X_3834_ _3834_/A vssd1 vssd1 vccd1 vccd1 _4504_/D sky130_fd_sc_hd__clkbuf_1
X_3765_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3765_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3696_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3696_/X sky130_fd_sc_hd__buf_2
X_2716_ _4357_/X _2713_/A _2317_/X _2715_/X vssd1 vssd1 vccd1 vccd1 _2716_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2647_ _4635_/Q vssd1 vssd1 vccd1 vccd1 _2703_/A sky130_fd_sc_hd__inv_2
XANTENNA__4342__A1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2578_ _4631_/Q vssd1 vssd1 vccd1 vccd1 _2721_/A sky130_fd_sc_hd__inv_2
XFILLER_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4317_ _4085_/X _4423_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4317_/X sky130_fd_sc_hd__mux2_1
X_4248_ _3992_/X _3989_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _4248_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4179_ _4146_/A _4146_/B _4147_/B vssd1 vssd1 vccd1 vccd1 _4180_/A sky130_fd_sc_hd__a21bo_1
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input49_A data_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3974__B _4250_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3550_ _4221_/X _4676_/Q _3554_/S vssd1 vssd1 vccd1 vccd1 _3551_/A sky130_fd_sc_hd__mux2_1
X_2501_ _4117_/A vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4324__A1 _4372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3481_ _3481_/A vssd1 vssd1 vccd1 vccd1 _4708_/D sky130_fd_sc_hd__clkbuf_1
X_2432_ _2317_/X _2319_/Y _2320_/Y vssd1 vssd1 vccd1 vccd1 _2433_/B sky130_fd_sc_hd__o21ai_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2886__A1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2363_ _3150_/A _2351_/B _2360_/X _2361_/X vssd1 vssd1 vccd1 vccd1 _2407_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4297__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4102_ _4102_/A vssd1 vssd1 vccd1 vccd1 _4102_/X sky130_fd_sc_hd__clkbuf_1
X_2294_ _4604_/Q _2293_/Y _2288_/B vssd1 vssd1 vccd1 vccd1 _2437_/B sky130_fd_sc_hd__o21ai_1
XFILLER_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4033_ _4036_/A _4033_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4033_/Y sky130_fd_sc_hd__nor3_1
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4045__B _4250_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3817_ _4514_/Q _3816_/X _4385_/X _3814_/X vssd1 vssd1 vccd1 vccd1 _4514_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3748_ _4563_/Q _3743_/X _2824_/A _3744_/X vssd1 vssd1 vccd1 vccd1 _4563_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4061__A _4109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3679_ _3717_/A vssd1 vssd1 vccd1 vccd1 _3696_/A sky130_fd_sc_hd__buf_4
Xoutput140 _3341_/A vssd1 vssd1 vccd1 vccd1 sb_hit sky130_fd_sc_hd__buf_2
XANTENNA__2877__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4410__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4701_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4401__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3817__B1 _4385_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2981_ _4443_/Q _2980_/Y _2998_/B vssd1 vssd1 vccd1 vccd1 _2991_/B sky130_fd_sc_hd__o21ai_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3985__A _3985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4720_ _4740_/CLK _4720_/D vssd1 vssd1 vccd1 vccd1 _4720_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_41_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4737_/CLK sky130_fd_sc_hd__clkbuf_16
X_4651_ _4742_/CLK _4651_/D vssd1 vssd1 vccd1 vccd1 _4651_/Q sky130_fd_sc_hd__dfxtp_1
Xinput20 addr_in[27] vssd1 vssd1 vccd1 vccd1 _2545_/A sky130_fd_sc_hd__buf_4
Xinput31 addr_in[8] vssd1 vssd1 vccd1 vccd1 _2472_/A sky130_fd_sc_hd__buf_6
X_3602_ _3602_/A vssd1 vssd1 vccd1 vccd1 _3602_/X sky130_fd_sc_hd__buf_2
Xinput53 data_in[28] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_4
Xinput42 data_in[18] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_2
X_4582_ _4583_/CLK _4582_/D vssd1 vssd1 vccd1 vccd1 _4582_/Q sky130_fd_sc_hd__dfxtp_1
Xinput64 data_in[9] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
X_3533_ _3533_/A vssd1 vssd1 vccd1 vccd1 _4684_/D sky130_fd_sc_hd__clkbuf_1
X_3464_ _4290_/X _4715_/Q _3464_/S vssd1 vssd1 vccd1 vccd1 _3465_/A sky130_fd_sc_hd__mux2_1
X_2415_ _2412_/X _2414_/X _2409_/X _2410_/Y vssd1 vssd1 vccd1 vccd1 _2415_/Y sky130_fd_sc_hd__a22oi_1
X_3395_ _3418_/S vssd1 vssd1 vccd1 vccd1 _3412_/S sky130_fd_sc_hd__buf_2
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2346_ _2344_/B _2343_/X _2344_/C vssd1 vssd1 vccd1 vccd1 _2346_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2277_ _4341_/X vssd1 vssd1 vccd1 vccd1 _2277_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4016_ _4020_/A _4035_/B _4017_/C vssd1 vssd1 vccd1 vccd1 _4016_/Y sky130_fd_sc_hd__nor3_1
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_32_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4746_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4395__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4565_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4386__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _4764_/Q vssd1 vssd1 vccd1 vccd1 _3287_/B sky130_fd_sc_hd__inv_2
X_3180_ _4547_/Q _3179_/Y _3076_/B vssd1 vssd1 vccd1 vccd1 _3181_/B sky130_fd_sc_hd__o21ai_1
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2964_ _3031_/A _2962_/Y _2963_/X vssd1 vssd1 vccd1 vccd1 _2964_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_14_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4556_/CLK sky130_fd_sc_hd__clkbuf_16
X_4703_ _4756_/CLK _4703_/D vssd1 vssd1 vccd1 vccd1 _4703_/Q sky130_fd_sc_hd__dfxtp_1
X_2895_ _2895_/A _2968_/A vssd1 vssd1 vccd1 vccd1 _2903_/C sky130_fd_sc_hd__or2_1
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2529__B1 _2543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4634_ _4634_/CLK _4634_/D vssd1 vssd1 vccd1 vccd1 _4634_/Q sky130_fd_sc_hd__dfxtp_1
X_4565_ _4565_/CLK _4565_/D vssd1 vssd1 vccd1 vccd1 _4565_/Q sky130_fd_sc_hd__dfxtp_1
X_3516_ _4272_/X _4691_/Q _3672_/S vssd1 vssd1 vccd1 vccd1 _3517_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4496_ _4629_/CLK _4496_/D vssd1 vssd1 vccd1 vccd1 _4496_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4377__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3447_ _3447_/A vssd1 vssd1 vccd1 vccd1 _4723_/D sky130_fd_sc_hd__clkbuf_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3378_ _4754_/Q _3373_/X _4241_/X _3375_/X vssd1 vssd1 vccd1 vccd1 _4754_/D sky130_fd_sc_hd__a22o_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _4595_/Q _2312_/Y _2336_/B vssd1 vssd1 vccd1 vccd1 _2329_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3257__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4368__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input31_A addr_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3799__A2 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2680_ _4647_/Q _2679_/Y _2676_/B vssd1 vssd1 vccd1 vccd1 _2792_/B sky130_fd_sc_hd__o21ai_1
X_4350_ _4181_/A _4146_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4350_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3301_ _3506_/A vssd1 vssd1 vccd1 vccd1 _3785_/A sky130_fd_sc_hd__inv_2
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ _4026_/Y input45/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4281_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4629_/CLK sky130_fd_sc_hd__clkbuf_16
X_3232_ _2456_/A _4559_/Q _2465_/A _4558_/Q vssd1 vssd1 vccd1 vccd1 _3260_/A sky130_fd_sc_hd__o22a_1
XFILLER_100_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3163_ _4192_/X _3175_/B vssd1 vssd1 vccd1 vccd1 _3163_/Y sky130_fd_sc_hd__nor2_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3094_ _3094_/A vssd1 vssd1 vccd1 vccd1 _3094_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3239__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3996_ _3996_/A vssd1 vssd1 vccd1 vccd1 _3996_/X sky130_fd_sc_hd__clkbuf_1
X_2947_ _2947_/A vssd1 vssd1 vccd1 vccd1 _2947_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4053__B _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2878_ _2878_/A _2878_/B _2878_/C _2878_/D vssd1 vssd1 vccd1 vccd1 _2878_/X sky130_fd_sc_hd__or4_1
X_4617_ _4751_/CLK _4617_/D vssd1 vssd1 vccd1 vccd1 _4617_/Q sky130_fd_sc_hd__dfxtp_1
X_4548_ _4583_/CLK _4548_/D vssd1 vssd1 vccd1 vccd1 _4548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4479_ _4757_/CLK _4479_/D vssd1 vssd1 vccd1 vccd1 _4479_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3650__B2 _3648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3323__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3850_ _4310_/X _4496_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3851_/A sky130_fd_sc_hd__mux2_1
X_2801_ _4470_/Q vssd1 vssd1 vccd1 vccd1 _2923_/A sky130_fd_sc_hd__inv_2
X_3781_ _3781_/A vssd1 vssd1 vccd1 vccd1 _4539_/D sky130_fd_sc_hd__clkbuf_1
X_2732_ _2353_/X _2727_/B _2779_/A _2731_/X vssd1 vssd1 vccd1 vccd1 _2781_/B sky130_fd_sc_hd__a22o_1
XANTENNA__3993__A _3993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2663_ _2668_/A _2660_/B _2661_/B vssd1 vssd1 vccd1 vccd1 _2663_/Y sky130_fd_sc_hd__a21boi_1
X_2594_ _2735_/A _2493_/A _2590_/Y _3380_/A vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__o22a_1
X_4402_ _4642_/Q _4599_/Q _4564_/Q _4464_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4402_/X sky130_fd_sc_hd__mux4_1
X_4333_ _4067_/X _4413_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4333_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4264_ _4263_/X input54/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4264_/X sky130_fd_sc_hd__mux2_2
XFILLER_99_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3215_ _4343_/X _3125_/Y _3214_/Y _3121_/Y _3124_/X vssd1 vssd1 vccd1 vccd1 _3216_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4195_ _3967_/Y _4042_/A _4195_/S vssd1 vssd1 vccd1 vccd1 _4195_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3146_ _3121_/Y _3129_/X _3216_/C _3144_/Y _3145_/Y vssd1 vssd1 vccd1 vccd1 _3146_/X
+ sky130_fd_sc_hd__o32a_1
X_3077_ _3234_/B _3198_/A _3196_/A _3196_/B vssd1 vssd1 vccd1 vccd1 _3152_/B sky130_fd_sc_hd__or4_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3979_ _4206_/X _3995_/B vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__and2_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3699__A1 _4595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3699__B2 _3697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4112__A2 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2222__A _4596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3000_ _4445_/Q _2998_/Y _2995_/B vssd1 vssd1 vccd1 vccd1 _3001_/B sky130_fd_sc_hd__o21ai_1
Xinput7 addr_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3500__B _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3902_ _4288_/X _4472_/Q _3958_/S vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__mux2_1
X_3833_ _4294_/X _4504_/Q _3841_/S vssd1 vssd1 vccd1 vccd1 _3834_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3764_ _3771_/A vssd1 vssd1 vccd1 vccd1 _3764_/X sky130_fd_sc_hd__clkbuf_2
X_3695_ _4597_/Q _3689_/X _2447_/A _3690_/X vssd1 vssd1 vccd1 vccd1 _4597_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2715_ _2702_/A _2702_/B _2703_/B vssd1 vssd1 vccd1 vccd1 _2715_/X sky130_fd_sc_hd__a21bo_1
X_2646_ _4636_/Q vssd1 vssd1 vccd1 vccd1 _2704_/A sky130_fd_sc_hd__inv_2
X_2577_ _2725_/A input4/X _2572_/X _2576_/X vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__o211a_1
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4316_ _4315_/X _4424_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4316_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4247_ _4246_/X _4375_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4247_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4059__A _4373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4178_ _4147_/A _4147_/B _4148_/B vssd1 vssd1 vccd1 vccd1 _4178_/X sky130_fd_sc_hd__a21bo_1
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3129_ _3124_/X _3214_/A _3216_/A vssd1 vssd1 vccd1 vccd1 _3129_/X sky130_fd_sc_hd__o21ba_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3837__S _3841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3844__A1 _4499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2500_ _2500_/A vssd1 vssd1 vccd1 vccd1 _4117_/A sky130_fd_sc_hd__inv_2
XFILLER_10_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3480_ _4225_/X _4708_/Q _3482_/S vssd1 vssd1 vccd1 vccd1 _3481_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2583__B2 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2431_ _2407_/A _2364_/X _2405_/X _2443_/C _2430_/X vssd1 vssd1 vccd1 vccd1 _2431_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2362_ _2360_/X _2361_/X _2353_/X _2356_/Y vssd1 vssd1 vccd1 vccd1 _2407_/B sky130_fd_sc_hd__o22ai_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2293_ _2293_/A _2293_/B vssd1 vssd1 vccd1 vccd1 _2293_/Y sky130_fd_sc_hd__nor2_1
X_4101_ _4430_/X _4103_/B vssd1 vssd1 vccd1 vccd1 _4102_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_4032_ _4036_/A _4032_/B _4036_/C vssd1 vssd1 vccd1 vccd1 _4032_/Y sky130_fd_sc_hd__nor3_1
XFILLER_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4260__A1 input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3816_ _3816_/A vssd1 vssd1 vccd1 vccd1 _3816_/X sky130_fd_sc_hd__clkbuf_4
X_3747_ _4564_/Q _3743_/X _2537_/A _3744_/X vssd1 vssd1 vccd1 vccd1 _4564_/D sky130_fd_sc_hd__a22o_1
X_3678_ _3678_/A _4770_/Q _3904_/C vssd1 vssd1 vccd1 vccd1 _3717_/A sky130_fd_sc_hd__or3_4
Xoutput130 _4478_/Q vssd1 vssd1 vccd1 vccd1 data_out[5] sky130_fd_sc_hd__buf_2
X_2629_ _4644_/Q vssd1 vssd1 vccd1 vccd1 _2667_/B sky130_fd_sc_hd__clkinv_2
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3762__B1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input61_A data_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2500__A _2500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3817__B2 _3814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2980_ _2980_/A _2980_/B vssd1 vssd1 vccd1 vccd1 _2980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4650_ _4737_/CLK _4650_/D vssd1 vssd1 vccd1 vccd1 _4650_/Q sky130_fd_sc_hd__dfxtp_1
Xinput21 addr_in[28] vssd1 vssd1 vccd1 vccd1 _2543_/A sky130_fd_sc_hd__buf_4
Xinput10 addr_in[18] vssd1 vssd1 vccd1 vccd1 _2464_/A sky130_fd_sc_hd__clkbuf_4
X_3601_ _3601_/A vssd1 vssd1 vccd1 vccd1 _3602_/A sky130_fd_sc_hd__inv_2
X_4581_ _4623_/CLK _4581_/D vssd1 vssd1 vccd1 vccd1 _4581_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3753__B1 _2452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput54 data_in[29] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_2
Xinput43 data_in[19] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_4
Xinput32 addr_in[9] vssd1 vssd1 vccd1 vccd1 _2474_/A sky130_fd_sc_hd__buf_6
Xinput65 hit_dtlb vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3532_ _4286_/X _4684_/Q _3536_/S vssd1 vssd1 vccd1 vccd1 _3533_/A sky130_fd_sc_hd__mux2_1
X_3463_ _3463_/A vssd1 vssd1 vccd1 vccd1 _4716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2414_ _2413_/A _2413_/B _2418_/B vssd1 vssd1 vccd1 vccd1 _2414_/X sky130_fd_sc_hd__a21bo_1
XFILLER_96_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3394_ _3569_/A _3576_/B _3594_/C vssd1 vssd1 vccd1 vccd1 _3418_/S sky130_fd_sc_hd__or3_4
X_2345_ _2345_/A vssd1 vssd1 vccd1 vccd1 _2345_/Y sky130_fd_sc_hd__inv_2
X_2276_ _2266_/X _2267_/X _2268_/X _2435_/A vssd1 vssd1 vccd1 vccd1 _2306_/B sky130_fd_sc_hd__o211ai_1
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3808__A1 _4520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4015_ _4039_/A vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4233__A1 _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4072__A _4094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2547__B2 _4602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4395__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3850__S _3852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2786__B2 _2798_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4386__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4215__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2963_ _4363_/X _2952_/X _4211_/X _2957_/Y vssd1 vssd1 vccd1 vccd1 _2963_/X sky130_fd_sc_hd__o22a_1
X_4702_ _4751_/CLK _4702_/D vssd1 vssd1 vccd1 vccd1 _4702_/Q sky130_fd_sc_hd__dfxtp_1
X_2894_ _2951_/A _2950_/A _2949_/A _4459_/Q vssd1 vssd1 vccd1 vccd1 _2938_/B sky130_fd_sc_hd__or4b_1
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2529__A1 _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _4634_/CLK _4633_/D vssd1 vssd1 vccd1 vccd1 _4633_/Q sky130_fd_sc_hd__dfxtp_1
X_4564_ _4642_/CLK _4564_/D vssd1 vssd1 vccd1 vccd1 _4564_/Q sky130_fd_sc_hd__dfxtp_2
X_3515_ _3515_/A vssd1 vssd1 vccd1 vccd1 _4692_/D sky130_fd_sc_hd__clkbuf_1
X_4495_ _4701_/CLK _4495_/D vssd1 vssd1 vccd1 vccd1 _4495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4377__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3446_ _4274_/X _4723_/Q _3728_/S vssd1 vssd1 vccd1 vccd1 _3447_/A sky130_fd_sc_hd__mux2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _4755_/Q _3373_/X _4237_/X _3375_/X vssd1 vssd1 vccd1 vccd1 _4755_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _2328_/A _2332_/B vssd1 vssd1 vccd1 vccd1 _2336_/B sky130_fd_sc_hd__or2_1
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2259_ _2272_/B _2259_/B vssd1 vssd1 vccd1 vccd1 _2259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4368__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input24_A addr_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3708__B1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2931__A1 _4470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3300_ _3965_/A _4195_/S vssd1 vssd1 vccd1 vccd1 _3506_/A sky130_fd_sc_hd__or2_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4280_ _4279_/X input46/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4280_/X sky130_fd_sc_hd__mux2_2
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _2466_/A _4558_/Q _2467_/A _4557_/Q vssd1 vssd1 vccd1 vccd1 _3263_/B sky130_fd_sc_hd__a22o_1
X_3162_ _4543_/Q _3161_/Y _3182_/B vssd1 vssd1 vccd1 vccd1 _3175_/B sky130_fd_sc_hd__o21ai_1
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3093_ _2266_/X _3086_/X _3087_/X _3217_/A vssd1 vssd1 vccd1 vccd1 _3115_/B sky130_fd_sc_hd__o211ai_1
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3947__B1 _2500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3995_ _4197_/X _3995_/B vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__and2_1
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2946_ _2944_/A _2944_/B _2944_/Y vssd1 vssd1 vccd1 vccd1 _2947_/A sky130_fd_sc_hd__a21oi_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2877_ input8/X _2949_/A _2876_/X vssd1 vssd1 vccd1 vccd1 _2878_/D sky130_fd_sc_hd__o21ai_1
X_4616_ _4760_/CLK _4616_/D vssd1 vssd1 vccd1 vccd1 _4616_/Q sky130_fd_sc_hd__dfxtp_1
X_4547_ _4583_/CLK _4547_/D vssd1 vssd1 vccd1 vccd1 _4547_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4478_ _4757_/CLK _4478_/D vssd1 vssd1 vccd1 vccd1 _4478_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3429_ _3429_/A vssd1 vssd1 vccd1 vccd1 _4731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3650__A2 _3647_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3938__B1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output130_A _4478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2800_ _2643_/Y _2800_/B vssd1 vssd1 vccd1 vccd1 _3969_/B sky130_fd_sc_hd__and2b_1
X_3780_ _4278_/X _4539_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3781_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_14_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2731_ _2725_/A _2725_/B _2725_/Y vssd1 vssd1 vccd1 vccd1 _2731_/X sky130_fd_sc_hd__a21o_1
X_2662_ _2667_/B _2661_/B _2661_/Y vssd1 vssd1 vccd1 vccd1 _2672_/A sky130_fd_sc_hd__a21oi_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4401_ _4641_/Q _4598_/Q _4563_/Q _4463_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4401_/X sky130_fd_sc_hd__mux4_1
X_2593_ _4620_/Q vssd1 vssd1 vccd1 vccd1 _2735_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_29_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4332_ _4331_/X _4417_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4332_/X sky130_fd_sc_hd__mux2_1
X_4263_ _4037_/Y input54/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4263_/X sky130_fd_sc_hd__mux2_1
X_3214_ _3214_/A vssd1 vssd1 vccd1 vccd1 _3214_/Y sky130_fd_sc_hd__inv_2
X_4194_ _4111_/X _3380_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4194_/X sky130_fd_sc_hd__mux2_4
XFILLER_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3145_ _3143_/B _3142_/X _3143_/C vssd1 vssd1 vccd1 vccd1 _3145_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3076_ _3076_/A _3076_/B vssd1 vssd1 vccd1 vccd1 _3196_/B sky130_fd_sc_hd__or2_1
XFILLER_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4064__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3978_ _4007_/B vssd1 vssd1 vccd1 vccd1 _3995_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2929_ _2926_/A _2926_/B _2926_/Y vssd1 vssd1 vccd1 vccd1 _2929_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3699__A2 _3696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4431__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 addr_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_6
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3901_ _3901_/A vssd1 vssd1 vccd1 vccd1 _4473_/D sky130_fd_sc_hd__clkbuf_1
X_3832_ _3900_/S vssd1 vssd1 vccd1 vccd1 _3841_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3763_ _4552_/Q _3757_/X input4/X _3758_/X vssd1 vssd1 vccd1 vccd1 _4552_/D sky130_fd_sc_hd__a22o_1
X_3694_ _4598_/Q _3689_/X _2824_/A _3690_/X vssd1 vssd1 vccd1 vccd1 _4598_/D sky130_fd_sc_hd__a22o_1
X_2714_ _4211_/X _2710_/Y _2711_/Y _2713_/Y vssd1 vssd1 vccd1 vccd1 _2788_/A sky130_fd_sc_hd__a22o_1
X_2645_ _2694_/A _2697_/A _2645_/C vssd1 vssd1 vccd1 vccd1 _2692_/A sky130_fd_sc_hd__or3_1
XFILLER_99_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4422__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4315_ _4087_/X _4424_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4315_/X sky130_fd_sc_hd__mux2_1
X_2576_ _2770_/A input2/X _2768_/A _2474_/A _2575_/X vssd1 vssd1 vccd1 vccd1 _2576_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4246_ _4044_/X _4375_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4246_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4059__B _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _4148_/A _4148_/B _4149_/B vssd1 vssd1 vccd1 vccd1 _4177_/X sky130_fd_sc_hd__a21bo_1
XFILLER_95_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3128_ _3121_/A _3121_/B _2321_/Y _3127_/Y vssd1 vssd1 vccd1 vccd1 _3216_/A sky130_fd_sc_hd__a22o_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ _4554_/Q vssd1 vssd1 vccd1 vccd1 _3148_/A sky130_fd_sc_hd__inv_2
XFILLER_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2592__A2 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4413__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2583__A2 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4404__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2430_ _2430_/A _2430_/B vssd1 vssd1 vccd1 vccd1 _2430_/X sky130_fd_sc_hd__or2_1
X_2361_ _2254_/A _2254_/B _2255_/B vssd1 vssd1 vccd1 vccd1 _2361_/X sky130_fd_sc_hd__a21bo_1
X_2292_ _2292_/A vssd1 vssd1 vccd1 vccd1 _2292_/X sky130_fd_sc_hd__clkbuf_2
X_4100_ _4100_/A vssd1 vssd1 vccd1 vccd1 _4100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4031_ _4039_/C vssd1 vssd1 vccd1 vccd1 _4036_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3815_ _4515_/Q _3809_/X _4386_/X _3814_/X vssd1 vssd1 vccd1 vccd1 _4515_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3746_ _4565_/Q _3743_/X _2816_/A _3744_/X vssd1 vssd1 vccd1 vccd1 _4565_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3677_ _4607_/Q _3601_/A _4262_/X _3602_/A vssd1 vssd1 vccd1 vccd1 _4607_/D sky130_fd_sc_hd__a22o_1
X_2628_ _4645_/Q vssd1 vssd1 vccd1 vccd1 _2667_/A sky130_fd_sc_hd__inv_2
Xoutput120 _4498_/Q vssd1 vssd1 vccd1 vccd1 data_out[25] sky130_fd_sc_hd__buf_2
Xoutput131 _4479_/Q vssd1 vssd1 vccd1 vccd1 data_out[6] sky130_fd_sc_hd__buf_2
X_2559_ _4640_/Q vssd1 vssd1 vccd1 vccd1 _2645_/C sky130_fd_sc_hd__inv_2
XFILLER_101_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4229_ _4228_/X input63/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4229_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2318__A _2318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3848__S _3852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input54_A data_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3817__A2 _3816_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ _4623_/CLK _4580_/D vssd1 vssd1 vccd1 vccd1 _4580_/Q sky130_fd_sc_hd__dfxtp_1
X_3600_ _3601_/A vssd1 vssd1 vccd1 vccd1 _3600_/X sky130_fd_sc_hd__buf_2
Xinput11 addr_in[19] vssd1 vssd1 vccd1 vccd1 _2455_/A sky130_fd_sc_hd__buf_4
Xinput22 addr_in[29] vssd1 vssd1 vccd1 vccd1 _2803_/A sky130_fd_sc_hd__buf_8
Xinput55 data_in[2] vssd1 vssd1 vccd1 vccd1 _3985_/A sky130_fd_sc_hd__buf_4
Xinput44 data_in[1] vssd1 vssd1 vccd1 vccd1 _3981_/A sky130_fd_sc_hd__buf_2
Xinput33 data_in[0] vssd1 vssd1 vccd1 vccd1 _3975_/A sky130_fd_sc_hd__clkbuf_2
X_3531_ _3531_/A vssd1 vssd1 vccd1 vccd1 _4685_/D sky130_fd_sc_hd__clkbuf_1
Xinput66 is_byte vssd1 vssd1 vccd1 vccd1 _4367_/S sky130_fd_sc_hd__buf_12
X_3462_ _4288_/X _4716_/Q _3464_/S vssd1 vssd1 vccd1 vccd1 _3463_/A sky130_fd_sc_hd__mux2_1
X_3393_ _3974_/A _3972_/A _4029_/C _3352_/A vssd1 vssd1 vccd1 vccd1 _3594_/C sky130_fd_sc_hd__o211a_1
X_2413_ _2413_/A _2413_/B vssd1 vssd1 vccd1 vccd1 _2418_/B sky130_fd_sc_hd__or2_1
XFILLER_97_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2344_ _2344_/A _2344_/B _2344_/C _2343_/X vssd1 vssd1 vccd1 vccd1 _2434_/A sky130_fd_sc_hd__or4b_1
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3269__B1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2275_ _3092_/A _2275_/B vssd1 vssd1 vccd1 vccd1 _2435_/A sky130_fd_sc_hd__or2_1
XANTENNA__3808__A2 _3802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4014_ _4014_/A vssd1 vssd1 vccd1 vccd1 _4039_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_3_0_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2547__A2 _4603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3729_ _3729_/A vssd1 vssd1 vccd1 vccd1 _4573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3432__A _3484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2511__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4202__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3342__A _3342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2962_ _4357_/X _2959_/A _2317_/A _2961_/X vssd1 vssd1 vccd1 vccd1 _2962_/Y sky130_fd_sc_hd__a22oi_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4701_/CLK _4701_/D vssd1 vssd1 vccd1 vccd1 _4701_/Q sky130_fd_sc_hd__dfxtp_1
X_4632_ _4634_/CLK _4632_/D vssd1 vssd1 vccd1 vccd1 _4632_/Q sky130_fd_sc_hd__dfxtp_2
X_2893_ _4457_/Q vssd1 vssd1 vccd1 vccd1 _2950_/A sky130_fd_sc_hd__inv_2
X_4563_ _4565_/CLK _4563_/D vssd1 vssd1 vccd1 vccd1 _4563_/Q sky130_fd_sc_hd__dfxtp_2
X_3514_ _4270_/X _4692_/Q _3514_/S vssd1 vssd1 vccd1 vccd1 _3515_/A sky130_fd_sc_hd__mux2_1
X_4494_ _4637_/CLK _4494_/D vssd1 vssd1 vccd1 vccd1 _4494_/Q sky130_fd_sc_hd__dfxtp_4
X_3445_ _3445_/A vssd1 vssd1 vccd1 vccd1 _4724_/D sky130_fd_sc_hd__clkbuf_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _4756_/Q _3373_/X _4233_/X _3375_/X vssd1 vssd1 vccd1 vccd1 _4756_/D sky130_fd_sc_hd__a22o_1
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _2327_/A vssd1 vssd1 vccd1 vccd1 _2327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2258_ _2273_/A _2258_/B vssd1 vssd1 vccd1 vccd1 _2259_/B sky130_fd_sc_hd__or2_1
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3662__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4083__A _4094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3861__S _3863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input17_A addr_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3653__B1 _2507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3337__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output85_A _4529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _2460_/A _4556_/Q _2462_/A _4557_/Q vssd1 vssd1 vccd1 vccd1 _3260_/B sky130_fd_sc_hd__o22a_1
X_3161_ _3161_/A _3161_/B vssd1 vssd1 vccd1 vccd1 _3161_/Y sky130_fd_sc_hd__nor2_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__A _4663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3092_ _3092_/A _3092_/B vssd1 vssd1 vccd1 vccd1 _3217_/A sky130_fd_sc_hd__or2_1
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3800__A _3814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3644__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3994_ _4036_/B _3994_/B vssd1 vssd1 vccd1 vccd1 _3994_/Y sky130_fd_sc_hd__nor2_1
X_2945_ _4461_/Q _2944_/Y _2941_/X vssd1 vssd1 vccd1 vccd1 _2945_/Y sky130_fd_sc_hd__o21ai_1
X_2876_ _2521_/A _4461_/Q _2453_/A _4460_/Q vssd1 vssd1 vccd1 vccd1 _2876_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4615_ _4755_/CLK _4615_/D vssd1 vssd1 vccd1 vccd1 _4615_/Q sky130_fd_sc_hd__dfxtp_1
X_4546_ _4621_/CLK _4546_/D vssd1 vssd1 vccd1 vccd1 _4546_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4477_ _4755_/CLK _4477_/D vssd1 vssd1 vccd1 vccd1 _4477_/Q sky130_fd_sc_hd__dfxtp_1
X_3428_ _4260_/X _4731_/Q _3430_/S vssd1 vssd1 vccd1 vccd1 _3429_/A sky130_fd_sc_hd__mux2_1
X_3359_ _3359_/A vssd1 vssd1 vccd1 vccd1 _4759_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input9_A addr_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3710__A _3717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3635__B1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4115__A1 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output123_A _4501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3620__A _3634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2730_ _4359_/X vssd1 vssd1 vccd1 vccd1 _2779_/A sky130_fd_sc_hd__inv_2
X_2661_ _2667_/B _2661_/B vssd1 vssd1 vccd1 vccd1 _2661_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3067__A _4547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4400_ _4640_/Q _4597_/Q _4562_/Q _4462_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4400_/X sky130_fd_sc_hd__mux4_1
XFILLER_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2592_ _2590_/Y _3380_/A _2591_/Y input1/X vssd1 vssd1 vccd1 vccd1 _2592_/X sky130_fd_sc_hd__a211o_1
X_4331_ _4069_/X _4417_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4331_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4262_ _4261_/X _3975_/A _4354_/S vssd1 vssd1 vccd1 vccd1 _4262_/X sky130_fd_sc_hd__mux2_2
X_3213_ _3208_/A _3160_/Y _3195_/X _3225_/C _3212_/X vssd1 vssd1 vccd1 vccd1 _3213_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4193_ _4123_/X _2506_/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4193_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4409__A2 _4571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3144_ _3144_/A vssd1 vssd1 vccd1 vccd1 _3144_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3075_ _3178_/A _3182_/A _3075_/C _3182_/B vssd1 vssd1 vccd1 vccd1 _3076_/B sky130_fd_sc_hd__or4_2
XFILLER_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3977_ _4032_/B _3994_/B vssd1 vssd1 vccd1 vccd1 _3977_/Y sky130_fd_sc_hd__nor2_1
X_2928_ _3035_/B vssd1 vssd1 vccd1 vccd1 _2928_/Y sky130_fd_sc_hd__inv_2
X_2859_ _4444_/Q vssd1 vssd1 vccd1 vccd1 _2998_/A sky130_fd_sc_hd__inv_2
XANTENNA__4345__A1 _4153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4529_ _4565_/CLK _4529_/D vssd1 vssd1 vccd1 vccd1 _4529_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4300__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3608__A0 _4284_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3586__S _3586_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4431__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4210__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3615__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput9 addr_in[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_4
X_3900_ _4252_/X _4473_/Q _3900_/S vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _3887_/A vssd1 vssd1 vccd1 vccd1 _3900_/S sky130_fd_sc_hd__buf_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3762_ _4553_/Q _3757_/X input5/X _3758_/X vssd1 vssd1 vccd1 vccd1 _4553_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3693_ _4599_/Q _3689_/X _2537_/A _3690_/X vssd1 vssd1 vccd1 vccd1 _4599_/D sky130_fd_sc_hd__a22o_1
X_2713_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2713_/Y sky130_fd_sc_hd__inv_2
X_2644_ _4638_/Q vssd1 vssd1 vccd1 vccd1 _2697_/A sky130_fd_sc_hd__inv_2
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2575_ _4626_/Q _2473_/X _4627_/Q _2513_/X vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4422__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4314_ _4313_/X _4425_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4314_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4245_ _4244_/X _3993_/A _4354_/S vssd1 vssd1 vccd1 vccd1 _4245_/X sky130_fd_sc_hd__mux2_2
X_4176_ _4149_/A _4149_/B _4150_/B vssd1 vssd1 vccd1 vccd1 _4176_/X sky130_fd_sc_hd__a21bo_1
XFILLER_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3127_ _3127_/A vssd1 vssd1 vccd1 vccd1 _3127_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ _4555_/Q vssd1 vssd1 vccd1 vccd1 _3060_/A sky130_fd_sc_hd__inv_2
XFILLER_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4075__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4413__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_13_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_28_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4205__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4404__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3345__A _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2360_ _3156_/A vssd1 vssd1 vccd1 vccd1 _2360_/X sky130_fd_sc_hd__clkbuf_2
X_2291_ _4347_/X vssd1 vssd1 vccd1 vccd1 _2292_/A sky130_fd_sc_hd__inv_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4030_ _4039_/A vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4690_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3814_ _3814_/A vssd1 vssd1 vccd1 vccd1 _3814_/X sky130_fd_sc_hd__clkbuf_4
X_3745_ _4566_/Q _3743_/X _2815_/A _3744_/X vssd1 vssd1 vccd1 vccd1 _4566_/D sky130_fd_sc_hd__a22o_1
Xoutput110 _4489_/Q vssd1 vssd1 vccd1 vccd1 data_out[16] sky130_fd_sc_hd__buf_2
X_3676_ _4608_/Q _3601_/A _4233_/X _3602_/A vssd1 vssd1 vccd1 vccd1 _4608_/D sky130_fd_sc_hd__a22o_1
Xoutput121 _4499_/Q vssd1 vssd1 vccd1 vccd1 data_out[26] sky130_fd_sc_hd__buf_2
Xoutput132 _4480_/Q vssd1 vssd1 vccd1 vccd1 data_out[7] sky130_fd_sc_hd__buf_2
X_2627_ _4649_/Q _2536_/X _4642_/Q _4153_/A _2626_/X vssd1 vssd1 vccd1 vccd1 _2637_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_99_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2558_ _4639_/Q vssd1 vssd1 vccd1 vccd1 _2694_/A sky130_fd_sc_hd__inv_2
X_2489_ _2489_/A _2489_/B _2489_/C _2489_/D vssd1 vssd1 vccd1 vccd1 _2489_/Y sky130_fd_sc_hd__nor4_1
X_4228_ _4011_/Y input63/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4228_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4159_ _4160_/B vssd1 vssd1 vccd1 vccd1 _4159_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_35_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4735_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4398__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input47_A data_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_26_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4600_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2244__A _4665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 addr_in[1] vssd1 vssd1 vccd1 vccd1 _3380_/A sky130_fd_sc_hd__buf_12
Xinput34 data_in[10] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_4
Xinput45 data_in[20] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 addr_in[2] vssd1 vssd1 vccd1 vccd1 _2493_/A sky130_fd_sc_hd__buf_6
X_3530_ _4284_/X _4685_/Q _3530_/S vssd1 vssd1 vccd1 vccd1 _3531_/A sky130_fd_sc_hd__mux2_1
Xinput67 reset vssd1 vssd1 vccd1 vccd1 _3965_/A sky130_fd_sc_hd__buf_6
Xinput56 data_in[30] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_2
XANTENNA__4389__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3461_ _3461_/A vssd1 vssd1 vccd1 vccd1 _4717_/D sky130_fd_sc_hd__clkbuf_1
X_2412_ _2412_/A vssd1 vssd1 vccd1 vccd1 _2412_/X sky130_fd_sc_hd__clkbuf_2
X_3392_ _3392_/A _3392_/B vssd1 vssd1 vccd1 vccd1 _4029_/C sky130_fd_sc_hd__or2_2
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2343_ _4210_/X _2337_/X _2340_/X _2341_/X vssd1 vssd1 vccd1 vccd1 _2343_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3269__A1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2274_ _4602_/Q _2259_/Y _2293_/B vssd1 vssd1 vccd1 vccd1 _2275_/B sky130_fd_sc_hd__o21ai_1
X_4013_ _4013_/A _4034_/B _4017_/C vssd1 vssd1 vccd1 vccd1 _4013_/Y sky130_fd_sc_hd__nor3_1
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_clk clkbuf_opt_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4695_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3728_ _4256_/X _4573_/Q _3728_/S vssd1 vssd1 vccd1 vccd1 _3729_/A sky130_fd_sc_hd__mux2_1
X_3659_ _4621_/Q _3654_/X _2492_/A _3655_/X vssd1 vssd1 vccd1 vccd1 _4621_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3432__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3859__S _3863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2961_ _2949_/A _2949_/B _2950_/B vssd1 vssd1 vccd1 vccd1 _2961_/X sky130_fd_sc_hd__a21bo_1
XFILLER_15_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4737_/CLK _4700_/D vssd1 vssd1 vccd1 vccd1 _4700_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4631_ _4634_/CLK _4631_/D vssd1 vssd1 vccd1 vccd1 _4631_/Q sky130_fd_sc_hd__dfxtp_2
X_2892_ _4458_/Q vssd1 vssd1 vccd1 vccd1 _2951_/A sky130_fd_sc_hd__inv_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4562_ _4565_/CLK _4562_/D vssd1 vssd1 vccd1 vccd1 _4562_/Q sky130_fd_sc_hd__dfxtp_2
X_3513_ _3513_/A vssd1 vssd1 vccd1 vccd1 _4693_/D sky130_fd_sc_hd__clkbuf_1
X_4493_ _4740_/CLK _4493_/D vssd1 vssd1 vccd1 vccd1 _4493_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3444_ _4272_/X _4724_/Q _3728_/S vssd1 vssd1 vccd1 vccd1 _3445_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_6_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4634_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _3375_/A vssd1 vssd1 vccd1 vccd1 _3375_/X sky130_fd_sc_hd__buf_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _4366_/X vssd1 vssd1 vccd1 vccd1 _2327_/A sky130_fd_sc_hd__inv_2
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2257_ _2273_/B _2273_/D vssd1 vssd1 vccd1 vccd1 _2258_/B sky130_fd_sc_hd__or2_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3662__B2 _3634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4303__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3653__B2 _3648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3618__A _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4213__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output78_A _4523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3154_/X _3156_/X _3208_/B _3208_/D vssd1 vssd1 vccd1 vccd1 _3160_/Y sky130_fd_sc_hd__a31oi_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3091_ _4567_/Q _3082_/Y _3105_/B vssd1 vssd1 vccd1 vccd1 _3092_/B sky130_fd_sc_hd__o21ai_1
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3993_ _3993_/A vssd1 vssd1 vccd1 vccd1 _4036_/B sky130_fd_sc_hd__clkinv_2
X_2944_ _2944_/A _2944_/B vssd1 vssd1 vccd1 vccd1 _2944_/Y sky130_fd_sc_hd__nor2_1
X_2875_ _4456_/Q vssd1 vssd1 vccd1 vccd1 _2949_/A sky130_fd_sc_hd__inv_2
X_4614_ _4760_/CLK _4614_/D vssd1 vssd1 vccd1 vccd1 _4614_/Q sky130_fd_sc_hd__dfxtp_1
X_4545_ _4621_/CLK _4545_/D vssd1 vssd1 vccd1 vccd1 _4545_/Q sky130_fd_sc_hd__dfxtp_2
X_4476_ _4757_/CLK _4476_/D vssd1 vssd1 vccd1 vccd1 _4476_/Q sky130_fd_sc_hd__dfxtp_4
X_3427_ _3427_/A vssd1 vssd1 vccd1 vccd1 _4732_/D sky130_fd_sc_hd__clkbuf_1
X_3358_ _4221_/X _4759_/Q _3420_/S vssd1 vssd1 vccd1 vccd1 _3359_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _2309_/A _2309_/B vssd1 vssd1 vccd1 vccd1 _2310_/B sky130_fd_sc_hd__or2_1
X_3289_ _3341_/A _3342_/A _3289_/C input65/X vssd1 vssd1 vccd1 vccd1 _3325_/B sky130_fd_sc_hd__or4b_4
XANTENNA__3635__A1 _4639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4094__A _4094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2610__A2 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3872__S _3874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3571__B1 _4665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3874__A1 _4485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output116_A _4494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2660_ _2668_/A _2660_/B vssd1 vssd1 vccd1 vccd1 _2661_/B sky130_fd_sc_hd__or2_1
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2591_ _4618_/Q vssd1 vssd1 vccd1 vccd1 _2591_/Y sky130_fd_sc_hd__inv_2
X_4330_ _4329_/X _4418_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4330_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4261_ _3980_/X _3975_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _4261_/X sky130_fd_sc_hd__mux2_1
X_3212_ _3212_/A _3212_/B vssd1 vssd1 vccd1 vccd1 _3212_/X sky130_fd_sc_hd__or2_1
X_4192_ _4115_/X _2492_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4192_/X sky130_fd_sc_hd__mux2_2
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4409__A3 _4471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3143_ _3143_/A _3143_/B _3143_/C _3142_/X vssd1 vssd1 vccd1 vccd1 _3216_/C sky130_fd_sc_hd__or4b_1
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3074_ _3074_/A _3161_/A _3161_/B vssd1 vssd1 vccd1 vccd1 _3182_/B sky130_fd_sc_hd__or3_1
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4290__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3976_ _4006_/B vssd1 vssd1 vccd1 vccd1 _3994_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2927_ _4469_/Q _2926_/Y _2923_/B vssd1 vssd1 vccd1 vccd1 _3035_/B sky130_fd_sc_hd__o21ai_2
XFILLER_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2858_ _2854_/X _2856_/X _2857_/X vssd1 vssd1 vccd1 vccd1 _2858_/X sky130_fd_sc_hd__a21bo_1
X_2789_ _2789_/A _2789_/B _2789_/C _2717_/X vssd1 vssd1 vccd1 vccd1 _2798_/D sky130_fd_sc_hd__or4b_2
X_4528_ _4638_/CLK _4528_/D vssd1 vssd1 vccd1 vccd1 _4528_/Q sky130_fd_sc_hd__dfxtp_1
X_4459_ _4558_/CLK _4459_/D vssd1 vssd1 vccd1 vccd1 _4459_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3350__B _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4272__A1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3830_ _3965_/A _3830_/B vssd1 vssd1 vccd1 vccd1 _3887_/A sky130_fd_sc_hd__or2_2
X_3761_ _4554_/Q _3757_/X input6/X _3758_/X vssd1 vssd1 vccd1 vccd1 _4554_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2712_ _2703_/A _2703_/B _2704_/B vssd1 vssd1 vccd1 vccd1 _2713_/A sky130_fd_sc_hd__a21bo_1
XFILLER_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3692_ _4600_/Q _3689_/X _2816_/A _3690_/X vssd1 vssd1 vccd1 vccd1 _4600_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2643_ _4650_/Q _2643_/B vssd1 vssd1 vccd1 vccd1 _2643_/Y sky130_fd_sc_hd__nand2_1
X_2574_ _4627_/Q vssd1 vssd1 vccd1 vccd1 _2768_/A sky130_fd_sc_hd__inv_2
X_4313_ _4089_/X _4425_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4313_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4244_ _3996_/X _3993_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _4244_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4175_ _4175_/A vssd1 vssd1 vccd1 vccd1 _4175_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_67_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3126_ _4350_/X _3123_/Y _4343_/X _3125_/Y vssd1 vssd1 vccd1 vccd1 _3214_/A sky130_fd_sc_hd__o22a_1
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3057_ _4552_/Q vssd1 vssd1 vccd1 vccd1 _3151_/A sky130_fd_sc_hd__inv_2
XANTENNA__4263__A1 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3774__B1 _2498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3959_ _3959_/A vssd1 vssd1 vccd1 vccd1 _4436_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2329__A1 _4595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4311__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3829__A1 _2204_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4254__A1 _3985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2530__A _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3626__A _3633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4221__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2290_ _3104_/A _2290_/B vssd1 vssd1 vccd1 vccd1 _2305_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4245__A1 _3993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3813_ _4516_/Q _3809_/X _4387_/X _3807_/X vssd1 vssd1 vccd1 vccd1 _4516_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3744_ _3751_/A vssd1 vssd1 vccd1 vccd1 _3744_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3756__B1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3675_ _4609_/Q _3601_/A _4258_/X _3602_/A vssd1 vssd1 vccd1 vccd1 _4609_/D sky130_fd_sc_hd__a22o_1
Xoutput100 _4514_/Q vssd1 vssd1 vccd1 vccd1 addr_out[7] sky130_fd_sc_hd__buf_2
X_2626_ _2676_/A _2532_/A _2625_/Y _2535_/A vssd1 vssd1 vccd1 vccd1 _2626_/X sky130_fd_sc_hd__a22o_1
Xoutput122 _4500_/Q vssd1 vssd1 vccd1 vccd1 data_out[27] sky130_fd_sc_hd__buf_2
Xoutput111 _4490_/Q vssd1 vssd1 vccd1 vccd1 data_out[17] sky130_fd_sc_hd__buf_2
Xoutput133 _4481_/Q vssd1 vssd1 vccd1 vccd1 data_out[8] sky130_fd_sc_hd__buf_2
X_2557_ _2440_/X _2443_/Y _2556_/Y vssd1 vssd1 vccd1 vccd1 _3969_/A sky130_fd_sc_hd__o21ba_1
X_2488_ _2507_/A _2250_/A _2472_/A _2251_/A _2487_/X vssd1 vssd1 vccd1 vccd1 _2489_/D
+ sky130_fd_sc_hd__o221ai_4
XFILLER_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4227_ _4226_/X _4368_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4227_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4158_ _4158_/A _4158_/B vssd1 vssd1 vccd1 vccd1 _4160_/B sky130_fd_sc_hd__or2_1
XFILLER_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4086__B _4092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3109_ _4570_/Q _3099_/Y _3102_/X vssd1 vssd1 vccd1 vccd1 _3110_/B sky130_fd_sc_hd__o21ai_1
X_4089_ _4089_/A vssd1 vssd1 vccd1 vccd1 _4089_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4306__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3747__B1 _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4398__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4216__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 addr_in[20] vssd1 vssd1 vccd1 vccd1 _2452_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3738__B1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput46 data_in[21] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_4
Xinput24 addr_in[30] vssd1 vssd1 vccd1 vccd1 _2532_/A sky130_fd_sc_hd__buf_6
Xinput35 data_in[11] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_4
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput68 sb_re vssd1 vssd1 vccd1 vccd1 _2204_/A sky130_fd_sc_hd__clkbuf_1
Xinput57 data_in[31] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_2
XANTENNA__4389__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3460_ _4286_/X _4717_/Q _3464_/S vssd1 vssd1 vccd1 vccd1 _3461_/A sky130_fd_sc_hd__mux2_1
X_2411_ _4364_/X vssd1 vssd1 vccd1 vccd1 _2412_/A sky130_fd_sc_hd__inv_2
X_3391_ _4748_/Q _3374_/A _4262_/X _3375_/A vssd1 vssd1 vccd1 vccd1 _4748_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3910__B1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2342_ _3134_/A _2334_/B _2340_/X _2341_/X vssd1 vssd1 vccd1 vccd1 _2344_/C sky130_fd_sc_hd__a22o_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2273_ _2273_/A _2273_/B _2273_/C _2273_/D vssd1 vssd1 vccd1 vccd1 _2293_/B sky130_fd_sc_hd__or4_2
X_4012_ _4013_/A _4033_/B _4017_/C vssd1 vssd1 vccd1 vccd1 _4012_/Y sky130_fd_sc_hd__nor3_1
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2477__B1 _2474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4218__A1 _4373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_12_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3727_ _3727_/A vssd1 vssd1 vccd1 vccd1 _4574_/D sky130_fd_sc_hd__clkbuf_1
X_3658_ _4622_/Q _3654_/X _2500_/A _3655_/X vssd1 vssd1 vccd1 vccd1 _4622_/D sky130_fd_sc_hd__a22o_1
X_3589_ _3960_/S vssd1 vssd1 vccd1 vccd1 _3952_/S sky130_fd_sc_hd__buf_2
X_2609_ _2722_/A input6/X _2589_/A _2608_/X _2587_/X vssd1 vssd1 vccd1 vccd1 _2609_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_27_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4209__A1 _3997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2960_ _4211_/X _2957_/Y _2711_/Y _2959_/Y vssd1 vssd1 vccd1 vccd1 _3031_/A sky130_fd_sc_hd__a22o_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2891_ _2941_/A _2944_/A _2891_/C vssd1 vssd1 vccd1 vccd1 _2939_/A sky130_fd_sc_hd__or3_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4630_ _4634_/CLK _4630_/D vssd1 vssd1 vccd1 vccd1 _4630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4561_ _4638_/CLK _4561_/D vssd1 vssd1 vccd1 vccd1 _4561_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2702__B _2702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3512_ _4268_/X _4693_/Q _3514_/S vssd1 vssd1 vccd1 vccd1 _3513_/A sky130_fd_sc_hd__mux2_1
X_4492_ _4558_/CLK _4492_/D vssd1 vssd1 vccd1 vccd1 _4492_/Q sky130_fd_sc_hd__dfxtp_2
X_3443_ _3443_/A vssd1 vssd1 vccd1 vccd1 _4725_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3814__A _3814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3374_/A vssd1 vssd1 vccd1 vccd1 _3375_/A sky130_fd_sc_hd__inv_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _2320_/Y _2433_/D _2433_/C vssd1 vssd1 vccd1 vccd1 _2325_/X sky130_fd_sc_hd__o21ba_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2256_ _2256_/A _2332_/A _2311_/B _2318_/A vssd1 vssd1 vccd1 vccd1 _2273_/D sky130_fd_sc_hd__or4_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3662__A2 _3633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4759_ _4759_/CLK _4759_/D vssd1 vssd1 vccd1 vccd1 _4759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3653__A2 _3647_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2861__B1 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2803__A _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3634__A _3634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3090_ _3090_/A _3090_/B _3090_/C _3090_/D vssd1 vssd1 vccd1 vccd1 _3105_/B sky130_fd_sc_hd__or4_2
XFILLER_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _3992_/A vssd1 vssd1 vccd1 vccd1 _3992_/X sky130_fd_sc_hd__clkbuf_1
X_2943_ _2953_/A _2953_/B _2340_/A _2942_/X vssd1 vssd1 vccd1 vccd1 _2956_/A sky130_fd_sc_hd__a22o_1
XFILLER_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2874_ _2874_/A _2874_/B vssd1 vssd1 vccd1 vccd1 _2878_/C sky130_fd_sc_hd__nand2_1
X_4613_ _4760_/CLK _4613_/D vssd1 vssd1 vccd1 vccd1 _4613_/Q sky130_fd_sc_hd__dfxtp_1
X_4544_ _4621_/CLK _4544_/D vssd1 vssd1 vccd1 vccd1 _4544_/Q sky130_fd_sc_hd__dfxtp_1
X_4475_ _4750_/CLK _4475_/D vssd1 vssd1 vccd1 vccd1 _4475_/Q sky130_fd_sc_hd__dfxtp_1
X_3426_ _4264_/X _4732_/Q _3430_/S vssd1 vssd1 vccd1 vccd1 _3427_/A sky130_fd_sc_hd__mux2_1
X_3357_ _3357_/A vssd1 vssd1 vccd1 vccd1 _4760_/D sky130_fd_sc_hd__clkbuf_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2308_/A _2318_/A vssd1 vssd1 vccd1 vccd1 _2309_/B sky130_fd_sc_hd__or2_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3288_ _3288_/A vssd1 vssd1 vccd1 vccd1 _3289_/C sky130_fd_sc_hd__clkbuf_4
X_2239_ _4581_/Q vssd1 vssd1 vccd1 vccd1 _2249_/A sky130_fd_sc_hd__inv_2
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4314__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3571__A1 _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input22_A addr_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output109_A _4488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4224__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4434__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2590_ _4619_/Q vssd1 vssd1 vccd1 vccd1 _2590_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4260_ _4259_/X input56/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4260_/X sky130_fd_sc_hd__mux2_1
X_4191_ _4165_/X _4156_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4191_/X sky130_fd_sc_hd__mux2_1
X_3211_ _3209_/C _3210_/Y _3204_/X vssd1 vssd1 vccd1 vccd1 _3212_/B sky130_fd_sc_hd__o21ai_1
XFILLER_67_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3142_ _3136_/Y _3138_/X _2340_/X _3140_/Y vssd1 vssd1 vccd1 vccd1 _3142_/X sky130_fd_sc_hd__o22a_1
X_3073_ _4541_/Q _4540_/Q _3072_/Y vssd1 vssd1 vccd1 vccd1 _3161_/B sky130_fd_sc_hd__o21ai_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2825__B1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3975_ _3975_/A vssd1 vssd1 vccd1 vccd1 _4032_/B sky130_fd_sc_hd__clkinv_2
X_2926_ _2926_/A _2926_/B vssd1 vssd1 vccd1 vccd1 _2926_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2443__A _2443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2857_ _4114_/A _4443_/Q _2494_/A _4442_/Q vssd1 vssd1 vccd1 vccd1 _2857_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4425__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2788_ _2788_/A _2788_/B vssd1 vssd1 vccd1 vccd1 _2789_/B sky130_fd_sc_hd__or2_1
X_4527_ _4558_/CLK _4527_/D vssd1 vssd1 vccd1 vccd1 _4527_/Q sky130_fd_sc_hd__dfxtp_1
X_4458_ _4558_/CLK _4458_/D vssd1 vssd1 vccd1 vccd1 _4458_/Q sky130_fd_sc_hd__dfxtp_2
X_3409_ _3409_/A vssd1 vssd1 vccd1 vccd1 _4741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4389_ _4629_/Q _4586_/Q _4551_/Q _4451_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4389_/X sky130_fd_sc_hd__mux4_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4309__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3792__B2 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3883__S _3885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4416__S0 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4219__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3760_ _4555_/Q _3757_/X input7/X _3758_/X vssd1 vssd1 vccd1 vccd1 _4555_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3783__B2 _3303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3783__A1 _4537_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2711_ _4357_/X vssd1 vssd1 vccd1 vccd1 _2711_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4407__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3691_ _4601_/Q _3689_/X _2815_/A _3690_/X vssd1 vssd1 vccd1 vccd1 _4601_/D sky130_fd_sc_hd__a22o_1
X_2642_ _2619_/X _2637_/X _2641_/X vssd1 vssd1 vccd1 vccd1 _2643_/B sky130_fd_sc_hd__o21bai_2
X_2573_ _4628_/Q vssd1 vssd1 vccd1 vccd1 _2770_/A sky130_fd_sc_hd__inv_2
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4312_ _4311_/X _4426_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4312_/X sky130_fd_sc_hd__mux2_4
XFILLER_87_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4243_ _4242_/X _4376_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4243_/X sky130_fd_sc_hd__mux2_1
X_4174_ _4174_/A vssd1 vssd1 vccd1 vccd1 _4175_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_28_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3125_ _3116_/A _3119_/A _3117_/B vssd1 vssd1 vccd1 vccd1 _3125_/Y sky130_fd_sc_hd__a21boi_1
X_3056_ _4553_/Q vssd1 vssd1 vccd1 vccd1 _3242_/B sky130_fd_sc_hd__inv_2
XFILLER_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2274__A1 _4602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3958_ _4276_/X _4436_/Q _3958_/S vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2577__A2 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2909_ _2914_/A _2906_/B _2907_/B vssd1 vssd1 vccd1 vccd1 _2909_/Y sky130_fd_sc_hd__a21boi_2
X_3889_ _3889_/A vssd1 vssd1 vccd1 vccd1 _4479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3732__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3907__A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3812_ _4517_/Q _3809_/X _4388_/X _3807_/X vssd1 vssd1 vccd1 vccd1 _4517_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3743_ _3750_/A vssd1 vssd1 vccd1 vccd1 _3743_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3674_ _4610_/Q _3600_/X _4254_/X _3602_/X vssd1 vssd1 vccd1 vccd1 _4610_/D sky130_fd_sc_hd__a22o_1
X_2625_ _4649_/Q vssd1 vssd1 vccd1 vccd1 _2625_/Y sky130_fd_sc_hd__inv_2
Xoutput101 _4515_/Q vssd1 vssd1 vccd1 vccd1 addr_out[8] sky130_fd_sc_hd__buf_2
Xoutput123 _4501_/Q vssd1 vssd1 vccd1 vccd1 data_out[28] sky130_fd_sc_hd__buf_2
Xoutput112 _4491_/Q vssd1 vssd1 vccd1 vccd1 data_out[18] sky130_fd_sc_hd__buf_2
Xoutput134 _4482_/Q vssd1 vssd1 vccd1 vccd1 data_out[9] sky130_fd_sc_hd__buf_2
X_2556_ _4763_/Q _2556_/B vssd1 vssd1 vccd1 vccd1 _2556_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2487_ input5/X _2487_/B vssd1 vssd1 vccd1 vccd1 _2487_/X sky130_fd_sc_hd__or2_2
XFILLER_101_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4226_ _4056_/X _4368_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__mux2_1
X_4157_ _4157_/A _4157_/B vssd1 vssd1 vccd1 vccd1 _4158_/B sky130_fd_sc_hd__or2_1
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3108_ _4351_/X _3219_/B _4346_/X _3107_/Y vssd1 vssd1 vccd1 vccd1 _3114_/B sky130_fd_sc_hd__o22ai_1
XFILLER_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3692__B1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4088_ _4425_/X _4092_/B vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__and2_1
X_3039_ _3039_/A _3039_/B _2992_/X _2991_/Y vssd1 vssd1 vccd1 vccd1 _3039_/X sky130_fd_sc_hd__or4bb_1
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2631__A _4642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4322__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2806__A _4471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3738__A1 _4571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput36 data_in[12] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_4
Xinput14 addr_in[21] vssd1 vssd1 vccd1 vccd1 _2520_/A sky130_fd_sc_hd__buf_8
Xinput25 addr_in[31] vssd1 vssd1 vccd1 vccd1 _2535_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__4232__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput69 sb_we vssd1 vssd1 vccd1 vccd1 _2205_/A sky130_fd_sc_hd__buf_2
Xinput58 data_in[3] vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__buf_6
XANTENNA__2961__A2 _2949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput47 data_in[22] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2410_ _4583_/Q _2399_/Y _2413_/B vssd1 vssd1 vccd1 vccd1 _2410_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3390_ _4749_/Q _3374_/A _4258_/X _3375_/A vssd1 vssd1 vccd1 vccd1 _4749_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3910__A1 _4471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2341_ _2224_/A _2336_/X _2332_/Y vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__a21o_1
X_2272_ _2272_/A _2272_/B vssd1 vssd1 vccd1 vccd1 _2273_/C sky130_fd_sc_hd__or2_1
XFILLER_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4011_ _4013_/A _4032_/B _4017_/C vssd1 vssd1 vccd1 vccd1 _4011_/Y sky130_fd_sc_hd__nor3_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2477__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3426__A0 _4264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3726_ _4286_/X _4574_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3727_/A sky130_fd_sc_hd__mux2_1
X_3657_ _4623_/Q _3654_/X _2498_/A _3655_/X vssd1 vssd1 vccd1 vccd1 _4623_/D sky130_fd_sc_hd__a22o_1
X_3588_ _4354_/X _4353_/X _3588_/C vssd1 vssd1 vccd1 vccd1 _3960_/S sky130_fd_sc_hd__or3_4
X_2608_ _2725_/A input4/X _2589_/B _2607_/Y _2572_/X vssd1 vssd1 vccd1 vccd1 _2608_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2539_ _2532_/A _2288_/A _2535_/A _2286_/Y vssd1 vssd1 vccd1 vccd1 _2539_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4097__B _4103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4209_ _3998_/Y _3997_/A _4209_/S vssd1 vssd1 vccd1 vccd1 _4209_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4317__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input52_A data_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3656__B1 _2505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4227__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2890_ _4460_/Q vssd1 vssd1 vccd1 vccd1 _2944_/A sky130_fd_sc_hd__inv_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2271__A _4602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4560_ _4638_/CLK _4560_/D vssd1 vssd1 vccd1 vccd1 _4560_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3511_ _3511_/A vssd1 vssd1 vccd1 vccd1 _4694_/D sky130_fd_sc_hd__clkbuf_1
X_4491_ _4558_/CLK _4491_/D vssd1 vssd1 vccd1 vccd1 _4491_/Q sky130_fd_sc_hd__dfxtp_1
X_3442_ _4270_/X _4725_/Q _3442_/S vssd1 vssd1 vccd1 vccd1 _3443_/A sky130_fd_sc_hd__mux2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2698__A1 _4639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3373_ _3374_/A vssd1 vssd1 vccd1 vccd1 _3373_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _3121_/A _2314_/B _2321_/Y _2322_/X vssd1 vssd1 vccd1 vccd1 _2433_/C sky130_fd_sc_hd__a22o_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3830__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2255_ _2255_/A _2255_/B vssd1 vssd1 vccd1 vccd1 _2318_/A sky130_fd_sc_hd__or2_2
XFILLER_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2870__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2622__B2 _2543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4758_ _4759_/CLK _4758_/D vssd1 vssd1 vccd1 vccd1 _4758_/Q sky130_fd_sc_hd__dfxtp_1
X_3709_ _4587_/Q _3703_/X input4/X _3704_/X vssd1 vssd1 vccd1 vccd1 _4587_/D sky130_fd_sc_hd__a22o_1
X_4689_ _4746_/CLK _4689_/D vssd1 vssd1 vccd1 vccd1 _4689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3638__B1 _2464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2861__A1 _2500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3915__A _3922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3629__B1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _4199_/X _3995_/B vssd1 vssd1 vccd1 vccd1 _3992_/A sky130_fd_sc_hd__and2_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_26_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2942_ _2891_/C _2941_/X _2939_/Y vssd1 vssd1 vccd1 vccd1 _2942_/X sky130_fd_sc_hd__a21o_1
XANTENNA__2604__B2 _2505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2873_ _2839_/X _2851_/Y _2868_/X _2872_/X vssd1 vssd1 vccd1 vccd1 _2873_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__4357__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4612_ _4751_/CLK _4612_/D vssd1 vssd1 vccd1 vccd1 _4612_/Q sky130_fd_sc_hd__dfxtp_1
X_4543_ _4621_/CLK _4543_/D vssd1 vssd1 vccd1 vccd1 _4543_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4474_ _4759_/CLK _4474_/D vssd1 vssd1 vccd1 vccd1 _4474_/Q sky130_fd_sc_hd__dfxtp_1
X_3425_ _3425_/A vssd1 vssd1 vccd1 vccd1 _4733_/D sky130_fd_sc_hd__clkbuf_1
X_3356_ _4217_/X _4760_/Q _3420_/S vssd1 vssd1 vccd1 vccd1 _3357_/A sky130_fd_sc_hd__mux2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2540__B1 _4153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _4363_/X vssd1 vssd1 vccd1 vccd1 _3121_/A sky130_fd_sc_hd__inv_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3287_/A _3287_/B _4766_/Q vssd1 vssd1 vccd1 vccd1 _3288_/A sky130_fd_sc_hd__and3_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ _4582_/Q vssd1 vssd1 vccd1 vccd1 _2250_/A sky130_fd_sc_hd__inv_2
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3735__A _3771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4330__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input15_A addr_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4339__A1 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4434__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4240__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output83_A _4527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3210_ _3210_/A _3210_/B vssd1 vssd1 vccd1 vccd1 _3210_/Y sky130_fd_sc_hd__nor2_1
X_4190_ _4189_/X _3964_/Y _4338_/S vssd1 vssd1 vccd1 vccd1 _4190_/X sky130_fd_sc_hd__mux2_8
X_3141_ _2340_/X _3140_/Y _3134_/A _3134_/B vssd1 vssd1 vccd1 vccd1 _3143_/C sky130_fd_sc_hd__a22o_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3380__A _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3072_ _4663_/Q vssd1 vssd1 vccd1 vccd1 _3072_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2825__A1 _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4370__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3974_ _3974_/A _4250_/S vssd1 vssd1 vccd1 vccd1 _4209_/S sky130_fd_sc_hd__nor2_4
X_2925_ _2925_/A _2925_/B vssd1 vssd1 vccd1 vccd1 _2936_/A sky130_fd_sc_hd__nor2_1
X_2856_ _2493_/A _2980_/A _3380_/A _2852_/Y vssd1 vssd1 vccd1 vccd1 _2856_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4425__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2787_ _2317_/X _2715_/X _2716_/Y vssd1 vssd1 vccd1 vccd1 _2788_/B sky130_fd_sc_hd__o21ai_1
X_4526_ _4638_/CLK _4526_/D vssd1 vssd1 vccd1 vccd1 _4526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4457_ _4558_/CLK _4457_/D vssd1 vssd1 vccd1 vccd1 _4457_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3408_ _4274_/X _4741_/Q _3408_/S vssd1 vssd1 vccd1 vccd1 _3409_/A sky130_fd_sc_hd__mux2_1
X_4388_ _4628_/Q _4585_/Q _4550_/Q _4450_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4388_/X sky130_fd_sc_hd__mux4_2
XANTENNA_input7_A addr_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _4353_/X vssd1 vssd1 vccd1 vccd1 _3365_/A sky130_fd_sc_hd__inv_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4325__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3792__A2 _3788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4416__S1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2504__B1 _2505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output121_A _4499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4235__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3783__A2 _3508_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2710_ _2704_/A _2704_/B _2704_/Y vssd1 vssd1 vccd1 vccd1 _2710_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4407__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3690_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3690_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2641_ _2625_/Y _2535_/A _2626_/X _2640_/X vssd1 vssd1 vccd1 vccd1 _2641_/X sky130_fd_sc_hd__o22a_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2572_ _2656_/A input3/X vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__or2_1
X_4311_ _4091_/X _4426_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4311_/X sky130_fd_sc_hd__mux2_1
X_4242_ _4046_/X _4376_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4242_/X sky130_fd_sc_hd__mux2_1
X_4173_ _4150_/A _4150_/B _4151_/B vssd1 vssd1 vccd1 vccd1 _4174_/A sky130_fd_sc_hd__a21bo_1
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3124_ _4211_/X _3127_/A _4350_/X _3123_/Y vssd1 vssd1 vccd1 vccd1 _3124_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3055_ _3116_/A _3118_/A _3117_/A _4559_/Q vssd1 vssd1 vccd1 vccd1 _3119_/B sky130_fd_sc_hd__or4b_1
Xclkbuf_leaf_47_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4756_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ _3957_/A vssd1 vssd1 vccd1 vccd1 _4437_/D sky130_fd_sc_hd__clkbuf_1
X_2908_ _2913_/B _2907_/B _2907_/Y vssd1 vssd1 vccd1 vccd1 _2918_/A sky130_fd_sc_hd__a21oi_2
X_3888_ _4227_/X _4479_/Q _3896_/S vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__mux2_1
X_2839_ input4/X _2971_/A _2834_/X _2838_/X vssd1 vssd1 vccd1 vccd1 _2839_/X sky130_fd_sc_hd__o211a_1
X_4509_ _4769_/CLK _4509_/D vssd1 vssd1 vccd1 vccd1 _4509_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_38_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4759_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4411__A0 _4700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3894__S _3896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3923__A _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_29_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4637_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4402__A0 _4642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3811_ _4518_/Q _3809_/X _4389_/X _3807_/X vssd1 vssd1 vccd1 vccd1 _4518_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3742_ _4567_/Q _3734_/X _2545_/A _3737_/X vssd1 vssd1 vccd1 vccd1 _4567_/D sky130_fd_sc_hd__a22o_1
X_3673_ _3673_/A vssd1 vssd1 vccd1 vccd1 _4611_/D sky130_fd_sc_hd__clkbuf_1
X_2624_ _4648_/Q vssd1 vssd1 vccd1 vccd1 _2676_/A sky130_fd_sc_hd__inv_2
Xoutput124 _4502_/Q vssd1 vssd1 vccd1 vccd1 data_out[29] sky130_fd_sc_hd__buf_2
Xoutput113 _4492_/Q vssd1 vssd1 vccd1 vccd1 data_out[19] sky130_fd_sc_hd__buf_2
Xoutput102 _4516_/Q vssd1 vssd1 vccd1 vccd1 addr_out[9] sky130_fd_sc_hd__buf_2
X_2555_ _2528_/X _2550_/X _2554_/X vssd1 vssd1 vccd1 vccd1 _2556_/B sky130_fd_sc_hd__o21bai_2
Xoutput135 _4769_/Q vssd1 vssd1 vccd1 vccd1 drain_out sky130_fd_sc_hd__buf_2
X_2486_ _4136_/A _4590_/Q _4136_/B _4589_/Q _2485_/X vssd1 vssd1 vccd1 vccd1 _2489_/C
+ sky130_fd_sc_hd__a221o_1
X_4225_ _4224_/X input64/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4225_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4156_ _4156_/A _4156_/B vssd1 vssd1 vccd1 vccd1 _4157_/B sky130_fd_sc_hd__or2_1
X_3107_ _3105_/A _3105_/B _3105_/Y vssd1 vssd1 vccd1 vccd1 _3107_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _4087_/A vssd1 vssd1 vccd1 vccd1 _4087_/X sky130_fd_sc_hd__clkbuf_1
X_3038_ _3032_/A _2966_/X _3029_/X _3041_/D _3037_/X vssd1 vssd1 vccd1 vccd1 _3042_/A
+ sky130_fd_sc_hd__o221ai_4
XFILLER_43_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3743__A _3750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_1_0_clk_A clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 addr_in[22] vssd1 vssd1 vccd1 vccd1 _2447_/A sky130_fd_sc_hd__buf_6
Xinput26 addr_in[3] vssd1 vssd1 vccd1 vccd1 _2492_/A sky130_fd_sc_hd__buf_8
Xinput37 data_in[13] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
Xinput59 data_in[4] vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__buf_2
Xinput48 data_in[23] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2340_ _2340_/A vssd1 vssd1 vccd1 vccd1 _2340_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2271_ _4602_/Q vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__inv_2
X_4010_ _4020_/C vssd1 vssd1 vccd1 vccd1 _4017_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3725_ _4575_/Q _3696_/A input1/X _3697_/A vssd1 vssd1 vccd1 vccd1 _4575_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_9_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4583_/CLK sky130_fd_sc_hd__clkbuf_16
X_3656_ _4624_/Q _3654_/X _2505_/A _3655_/X vssd1 vssd1 vccd1 vccd1 _4624_/D sky130_fd_sc_hd__a22o_1
X_3587_ _3587_/A vssd1 vssd1 vccd1 vccd1 _4659_/D sky130_fd_sc_hd__clkbuf_1
X_2607_ _4628_/Q _2512_/X _4627_/Q _2513_/X _2575_/X vssd1 vssd1 vccd1 vccd1 _2607_/Y
+ sky130_fd_sc_hd__a221oi_2
XFILLER_88_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2538_ _2538_/A vssd1 vssd1 vccd1 vccd1 _4153_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4208_ _4002_/Y _4001_/A _4209_/S vssd1 vssd1 vccd1 vccd1 _4208_/X sky130_fd_sc_hd__mux2_1
X_2469_ _2457_/A _4594_/Q _2466_/A _4593_/Q vssd1 vssd1 vccd1 vccd1 _2519_/A sky130_fd_sc_hd__o22a_1
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3502__S _3514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4139_ _4134_/A _4134_/B _4136_/C vssd1 vssd1 vccd1 vccd1 _4139_/X sky130_fd_sc_hd__a21bo_1
XFILLER_56_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4333__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4393__A2 _4555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input45_A data_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4243__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3648__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3592__A0 _4256_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3510_ _4266_/X _4694_/Q _3514_/S vssd1 vssd1 vccd1 vccd1 _3511_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4490_ _4737_/CLK _4490_/D vssd1 vssd1 vccd1 vccd1 _4490_/Q sky130_fd_sc_hd__dfxtp_4
X_3441_ _3441_/A vssd1 vssd1 vccd1 vccd1 _4726_/D sky130_fd_sc_hd__clkbuf_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3372_/A vssd1 vssd1 vccd1 vccd1 _3374_/A sky130_fd_sc_hd__buf_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2321_/Y _2322_/X _4357_/X _2315_/X vssd1 vssd1 vccd1 vccd1 _2433_/D sky130_fd_sc_hd__o22ai_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _2254_/A _2254_/B vssd1 vssd1 vccd1 vccd1 _2255_/B sky130_fd_sc_hd__or2_1
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2622__A2 _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4757_ _4757_/CLK _4757_/D vssd1 vssd1 vccd1 vccd1 _4757_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3583__B1 _4661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3708_ _4588_/Q _3703_/X input5/X _3704_/X vssd1 vssd1 vccd1 vccd1 _4588_/D sky130_fd_sc_hd__a22o_1
X_4688_ _4746_/CLK _4688_/D vssd1 vssd1 vccd1 vccd1 _4688_/Q sky130_fd_sc_hd__dfxtp_1
X_3639_ _4635_/Q _3633_/X input9/X _3634_/X vssd1 vssd1 vccd1 vccd1 _4635_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4328__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3810__A1 _4519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4238__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3990_ _4035_/B _3994_/B vssd1 vssd1 vccd1 vccd1 _3990_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2604__A2 _2498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2941_ _2941_/A _2944_/A _2944_/B vssd1 vssd1 vccd1 vccd1 _2941_/X sky130_fd_sc_hd__or3_1
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3801__A1 _4525_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3801__B2 _3800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2872_ input7/X _2895_/A _2845_/X _2871_/X vssd1 vssd1 vccd1 vccd1 _2872_/X sky130_fd_sc_hd__o22a_1
X_4611_ _4744_/CLK _4611_/D vssd1 vssd1 vccd1 vccd1 _4611_/Q sky130_fd_sc_hd__dfxtp_1
X_4542_ _4621_/CLK _4542_/D vssd1 vssd1 vccd1 vccd1 _4542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4473_ _4701_/CLK _4473_/D vssd1 vssd1 vccd1 vccd1 _4473_/Q sky130_fd_sc_hd__dfxtp_1
X_3424_ _4213_/X _4733_/Q _3586_/S vssd1 vssd1 vccd1 vccd1 _3425_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3868__A1 _4488_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3355_ _3586_/S vssd1 vssd1 vccd1 vccd1 _3420_/S sky130_fd_sc_hd__buf_2
XANTENNA__3332__A3 _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2540__B2 _4599_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2540__A1 _2536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2306_ _2306_/A _2306_/B _2306_/C _2306_/D vssd1 vssd1 vccd1 vccd1 _2434_/C sky130_fd_sc_hd__or4_1
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3286_ _3286_/A vssd1 vssd1 vccd1 vccd1 _3341_/A sky130_fd_sc_hd__clkbuf_4
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _4583_/Q vssd1 vssd1 vccd1 vccd1 _2251_/A sky130_fd_sc_hd__inv_2
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3859__A1 _4492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3751__A _3751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4284__A1 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output76_A _4521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3140_ _4562_/Q _3137_/Y _3132_/X vssd1 vssd1 vccd1 vccd1 _3140_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2522__B2 _4595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3071_ _4542_/Q vssd1 vssd1 vccd1 vccd1 _3161_/A sky130_fd_sc_hd__inv_2
XANTENNA__4370__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4250_/S sky130_fd_sc_hd__clkbuf_4
X_2924_ _4470_/Q _2922_/Y _4471_/Q _2806_/Y _2923_/X vssd1 vssd1 vccd1 vccd1 _2925_/B
+ sky130_fd_sc_hd__a32o_1
X_2855_ _4442_/Q vssd1 vssd1 vccd1 vccd1 _2980_/A sky130_fd_sc_hd__inv_2
XFILLER_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2786_ _2781_/A _2734_/Y _2767_/X _2798_/C _2785_/X vssd1 vssd1 vccd1 vccd1 _2786_/X
+ sky130_fd_sc_hd__o221a_1
X_4525_ _4738_/CLK _4525_/D vssd1 vssd1 vccd1 vccd1 _4525_/Q sky130_fd_sc_hd__dfxtp_2
X_4456_ _4518_/CLK _4456_/D vssd1 vssd1 vccd1 vccd1 _4456_/Q sky130_fd_sc_hd__dfxtp_2
X_4387_ _4627_/Q _4584_/Q _4549_/Q _4449_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4387_/X sky130_fd_sc_hd__mux4_2
X_3407_ _3407_/A vssd1 vssd1 vccd1 vccd1 _4742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3338_ _3364_/A vssd1 vssd1 vccd1 vccd1 _3569_/A sky130_fd_sc_hd__clkbuf_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _2532_/A _3102_/A _2535_/A _3100_/Y vssd1 vssd1 vccd1 vccd1 _3269_/X sky130_fd_sc_hd__a22o_1
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4266__A1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3510__S _3514_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3777__B1 _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3241__A2 _4555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4341__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2504__A1 _2498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_25_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3701__B1 _2464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4257__A1 _3981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3768__B1 _2474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2640_ _2637_/A _2639_/X _2637_/B vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__4251__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2571_ _4629_/Q vssd1 vssd1 vccd1 vccd1 _2656_/A sky130_fd_sc_hd__inv_2
XANTENNA__3940__B1 _2474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4310_ _4309_/X _4427_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4310_/X sky130_fd_sc_hd__mux2_4
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4241_ _4240_/X _3997_/A _4354_/S vssd1 vssd1 vccd1 vccd1 _4241_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4172_ _4151_/A _4151_/B _4152_/B vssd1 vssd1 vccd1 vccd1 _4172_/X sky130_fd_sc_hd__a21bo_1
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4248__A1 _3989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3123_ _3117_/A _3117_/B _3118_/B vssd1 vssd1 vccd1 vccd1 _3123_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_82_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3054_ _4557_/Q vssd1 vssd1 vccd1 vccd1 _3117_/A sky130_fd_sc_hd__inv_2
XFILLER_70_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3759__B1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3956_ _4268_/X _4437_/Q _3960_/S vssd1 vssd1 vccd1 vccd1 _3957_/A sky130_fd_sc_hd__mux2_1
X_2907_ _2913_/B _2907_/B vssd1 vssd1 vccd1 vccd1 _2907_/Y sky130_fd_sc_hd__nor2_1
X_3887_ _3887_/A vssd1 vssd1 vccd1 vccd1 _3896_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2838_ input2/X _3014_/A _2474_/A _3012_/A _2837_/X vssd1 vssd1 vccd1 vccd1 _2838_/X
+ sky130_fd_sc_hd__o221a_1
X_2769_ _2768_/A _2768_/B _2770_/B vssd1 vssd1 vccd1 vccd1 _2769_/X sky130_fd_sc_hd__a21bo_1
X_4508_ _4618_/CLK _4508_/D vssd1 vssd1 vccd1 vccd1 _4508_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3931__B1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4439_ _4752_/CLK _4439_/D vssd1 vssd1 vccd1 vccd1 _4439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4336__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4411__A1 _4665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4246__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3810_ _4519_/Q _3809_/X _4390_/X _3807_/X vssd1 vssd1 vccd1 vccd1 _4519_/D sky130_fd_sc_hd__a22o_1
X_3741_ _4568_/Q _3734_/X _2543_/A _3737_/X vssd1 vssd1 vccd1 vccd1 _4568_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4402__A1 _4599_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3672_ _4256_/X _4611_/Q _3672_/S vssd1 vssd1 vccd1 vccd1 _3673_/A sky130_fd_sc_hd__mux2_1
X_2623_ _4647_/Q _4158_/A _4648_/Q _4160_/A vssd1 vssd1 vccd1 vccd1 _2637_/B sky130_fd_sc_hd__a22o_1
XANTENNA__3913__B1 _2543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2554_ _2535_/A _2286_/Y _2539_/X _2553_/X vssd1 vssd1 vccd1 vccd1 _2554_/X sky130_fd_sc_hd__o22a_1
Xoutput125 _4475_/Q vssd1 vssd1 vccd1 vccd1 data_out[2] sky130_fd_sc_hd__buf_2
Xoutput103 _4473_/Q vssd1 vssd1 vccd1 vccd1 data_out[0] sky130_fd_sc_hd__buf_2
Xoutput114 _4474_/Q vssd1 vssd1 vccd1 vccd1 data_out[1] sky130_fd_sc_hd__buf_2
Xoutput136 _2207_/B vssd1 vssd1 vccd1 vccd1 empty_out sky130_fd_sc_hd__buf_2
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2485_ input7/X _2255_/A input6/X _2254_/A vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4224_ _4012_/Y input64/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4224_/X sky130_fd_sc_hd__mux2_1
X_4155_ _4155_/A _4155_/B vssd1 vssd1 vccd1 vccd1 _4156_/B sky130_fd_sc_hd__or2_1
X_3106_ _4569_/Q _3105_/Y _3102_/B vssd1 vssd1 vccd1 vccd1 _3219_/B sky130_fd_sc_hd__o21a_1
XFILLER_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ _4424_/X _4092_/B vssd1 vssd1 vccd1 vccd1 _4087_/A sky130_fd_sc_hd__and2_1
XFILLER_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3037_ _3033_/Y _3034_/X _2937_/D _2936_/A _3036_/Y vssd1 vssd1 vccd1 vccd1 _3037_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3939_ _4450_/Q _3936_/X input2/X _3937_/X vssd1 vssd1 vccd1 vccd1 _4450_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2375__A _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput27 addr_in[4] vssd1 vssd1 vccd1 vccd1 _2500_/A sky130_fd_sc_hd__buf_6
Xinput16 addr_in[23] vssd1 vssd1 vccd1 vccd1 _2824_/A sky130_fd_sc_hd__buf_8
Xinput49 data_in[24] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_4
Xinput38 data_in[14] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2270_ _2916_/A vssd1 vssd1 vccd1 vccd1 _3092_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4773_ _4773_/CLK _4773_/D vssd1 vssd1 vccd1 vccd1 _4773_/Q sky130_fd_sc_hd__dfxtp_1
X_3724_ _4576_/Q _3696_/A _3380_/A _3697_/A vssd1 vssd1 vccd1 vccd1 _4576_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4005__A _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3655_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3655_/X sky130_fd_sc_hd__clkbuf_2
X_2606_ _2601_/X _2604_/X _2605_/X vssd1 vssd1 vccd1 vccd1 _2606_/X sky130_fd_sc_hd__a21bo_2
X_3586_ _4215_/X _4659_/Q _3586_/S vssd1 vssd1 vccd1 vccd1 _3587_/A sky130_fd_sc_hd__mux2_1
X_2537_ _2537_/A vssd1 vssd1 vccd1 vccd1 _2538_/A sky130_fd_sc_hd__inv_2
XFILLER_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2468_ _4147_/A _4593_/Q _4146_/A _4592_/Q vssd1 vssd1 vccd1 vccd1 _2524_/B sky130_fd_sc_hd__a22o_1
X_4207_ _4006_/Y _4005_/A _4209_/S vssd1 vssd1 vccd1 vccd1 _4207_/X sky130_fd_sc_hd__mux2_1
X_2399_ _2399_/A vssd1 vssd1 vccd1 vccd1 _2399_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4138_ _4136_/B _4136_/C _4135_/Y vssd1 vssd1 vccd1 vccd1 _4138_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4069_ _4069_/A vssd1 vssd1 vccd1 vccd1 _4069_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input38_A data_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3929__A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3440_ _4268_/X _4726_/Q _3442_/S vssd1 vssd1 vccd1 vccd1 _3441_/A sky130_fd_sc_hd__mux2_1
X_3371_ _3484_/A _3556_/B _3598_/C vssd1 vssd1 vccd1 vccd1 _3372_/A sky130_fd_sc_hd__or3_1
XFILLER_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2322_ _2310_/A _2310_/B _2310_/X vssd1 vssd1 vccd1 vccd1 _2322_/X sky130_fd_sc_hd__a21bo_1
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ _2487_/B _2354_/A _2355_/B vssd1 vssd1 vccd1 vccd1 _2254_/B sky130_fd_sc_hd__or3_1
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4756_ _4756_/CLK _4756_/D vssd1 vssd1 vccd1 vccd1 _4756_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3583__A1 _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3707_ _4589_/Q _3703_/X input6/X _3704_/X vssd1 vssd1 vccd1 vccd1 _4589_/D sky130_fd_sc_hd__a22o_1
X_4687_ _4740_/CLK _4687_/D vssd1 vssd1 vccd1 vccd1 _4687_/Q sky130_fd_sc_hd__dfxtp_1
X_3638_ _4636_/Q _3633_/X _2464_/A _3634_/X vssd1 vssd1 vccd1 vccd1 _4636_/D sky130_fd_sc_hd__a22o_1
X_3569_ _3569_/A _4353_/X _3581_/C vssd1 vssd1 vccd1 vccd1 _3570_/A sky130_fd_sc_hd__or3_1
XFILLER_29_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3271__B1 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4344__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3484__A _3484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2940_ _4463_/Q _2939_/Y _2914_/D vssd1 vssd1 vccd1 vccd1 _2953_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__4254__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2871_ input6/X _2968_/A _2851_/A _2870_/X _2849_/X vssd1 vssd1 vccd1 vccd1 _2871_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3801__A2 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4610_ _4706_/CLK _4610_/D vssd1 vssd1 vccd1 vccd1 _4610_/Q sky130_fd_sc_hd__dfxtp_1
X_4541_ _4695_/CLK _4541_/D vssd1 vssd1 vccd1 vccd1 _4541_/Q sky130_fd_sc_hd__dfxtp_1
X_4472_ _4737_/CLK _4472_/D vssd1 vssd1 vccd1 vccd1 _4472_/Q sky130_fd_sc_hd__dfxtp_1
X_3423_ _3423_/A vssd1 vssd1 vccd1 vccd1 _4734_/D sky130_fd_sc_hd__clkbuf_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3354_ _3569_/A _3576_/B _3572_/C vssd1 vssd1 vccd1 vccd1 _3586_/S sky130_fd_sc_hd__or3_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2305_/A _2305_/B _2305_/C _2305_/D vssd1 vssd1 vccd1 vccd1 _2306_/D sky130_fd_sc_hd__or4_1
XANTENNA__2738__A _4700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3285_ _3969_/A _3969_/B _3284_/X vssd1 vssd1 vccd1 vccd1 _3286_/A sky130_fd_sc_hd__or3b_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _4584_/Q vssd1 vssd1 vccd1 vccd1 _2413_/A sky130_fd_sc_hd__inv_2
XFILLER_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4428__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4739_ _4740_/CLK _4739_/D vssd1 vssd1 vccd1 vccd1 _4739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4339__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4419__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3011__A3 _3041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2558__A _4639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2522__A2 _4596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4249__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3070_ _4543_/Q vssd1 vssd1 vccd1 vccd1 _3074_/A sky130_fd_sc_hd__inv_2
XFILLER_85_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3972_ _3972_/A vssd1 vssd1 vccd1 vccd1 _4094_/A sky130_fd_sc_hd__buf_2
X_2923_ _2923_/A _2923_/B vssd1 vssd1 vccd1 vccd1 _2923_/X sky130_fd_sc_hd__or2_1
X_2854_ _3380_/A _2852_/Y input1/X _2853_/Y vssd1 vssd1 vccd1 vccd1 _2854_/X sky130_fd_sc_hd__a211o_1
XFILLER_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2785_ _2785_/A _2785_/B vssd1 vssd1 vccd1 vccd1 _2785_/X sky130_fd_sc_hd__or2_1
XANTENNA__4013__A _4013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4524_ _4737_/CLK _4524_/D vssd1 vssd1 vccd1 vccd1 _4524_/Q sky130_fd_sc_hd__dfxtp_2
X_4455_ _4589_/CLK _4455_/D vssd1 vssd1 vccd1 vccd1 _4455_/Q sky130_fd_sc_hd__dfxtp_2
X_4386_ _4626_/Q _4583_/Q _4548_/Q _4448_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4386_/X sky130_fd_sc_hd__mux4_2
X_3406_ _4272_/X _4742_/Q _3408_/S vssd1 vssd1 vccd1 vccd1 _3407_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3337_ _4354_/X vssd1 vssd1 vccd1 vccd1 _3364_/A sky130_fd_sc_hd__inv_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _2531_/A _4569_/Q _4160_/A _4570_/Q vssd1 vssd1 vccd1 vccd1 _3276_/B sky130_fd_sc_hd__a22o_1
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _4599_/Q vssd1 vssd1 vccd1 vccd1 _2273_/B sky130_fd_sc_hd__inv_2
X_3199_ _3198_/A _3198_/B _3198_/X vssd1 vssd1 vccd1 vccd1 _3199_/X sky130_fd_sc_hd__a21bo_1
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3226__B1 _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3701__B2 _3697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input20_A addr_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3937__A _3944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2570_ _2721_/B vssd1 vssd1 vccd1 vccd1 _2725_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4240_ _4000_/X _3997_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _4240_/X sky130_fd_sc_hd__mux2_1
X_4171_ _4152_/A _4152_/B _4153_/B vssd1 vssd1 vccd1 vccd1 _4171_/X sky130_fd_sc_hd__a21bo_1
X_3122_ _3118_/A _3118_/B _3118_/Y vssd1 vssd1 vccd1 vccd1 _3127_/A sky130_fd_sc_hd__a21oi_1
XFILLER_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3053_ _4558_/Q vssd1 vssd1 vccd1 vccd1 _3118_/A sky130_fd_sc_hd__inv_2
XFILLER_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3759__A1 _4556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3955_ _3955_/A vssd1 vssd1 vccd1 vccd1 _4438_/D sky130_fd_sc_hd__clkbuf_1
X_2906_ _2914_/A _2906_/B vssd1 vssd1 vccd1 vccd1 _2907_/B sky130_fd_sc_hd__or2_1
X_3886_ _3886_/A vssd1 vssd1 vccd1 vccd1 _4480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2837_ _2473_/X _4448_/Q _4130_/A _4449_/Q vssd1 vssd1 vccd1 vccd1 _2837_/X sky130_fd_sc_hd__o22a_1
X_2768_ _2768_/A _2768_/B vssd1 vssd1 vccd1 vccd1 _2770_/B sky130_fd_sc_hd__or2_1
X_4507_ _4618_/CLK _4507_/D vssd1 vssd1 vccd1 vccd1 _4507_/Q sky130_fd_sc_hd__dfxtp_4
X_2699_ _2697_/A _2697_/B _2697_/Y vssd1 vssd1 vccd1 vccd1 _2700_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__3931__A1 _4456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4438_ _4690_/CLK _4438_/D vssd1 vssd1 vccd1 vccd1 _4438_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3695__B1 _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4369_ _4741_/Q _4723_/Q _4690_/Q _4438_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4369_/X sky130_fd_sc_hd__mux4_2
XFILLER_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4411__A2 _4663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4352__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3757__A _3771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input68_A sb_re vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3686__B1 _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3438__A0 _4266_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3740_ _4569_/Q _3734_/X _2803_/A _3737_/X vssd1 vssd1 vccd1 vccd1 _4569_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4262__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3671_ _4612_/Q _3600_/X _4249_/X _3602_/X vssd1 vssd1 vccd1 vccd1 _4612_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2622_ _2674_/A _2803_/A _2679_/A _2543_/A vssd1 vssd1 vccd1 vccd1 _2637_/A sky130_fd_sc_hd__a22o_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput115 _4493_/Q vssd1 vssd1 vccd1 vccd1 data_out[20] sky130_fd_sc_hd__buf_2
X_2553_ _2550_/A _2552_/X _2550_/B vssd1 vssd1 vccd1 vccd1 _2553_/X sky130_fd_sc_hd__o21ba_1
Xoutput104 _4483_/Q vssd1 vssd1 vccd1 vccd1 data_out[10] sky130_fd_sc_hd__buf_2
Xoutput137 _3289_/C vssd1 vssd1 vccd1 vccd1 full_out sky130_fd_sc_hd__buf_2
XANTENNA__3606__S _3606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput126 _4503_/Q vssd1 vssd1 vccd1 vccd1 data_out[30] sky130_fd_sc_hd__buf_2
X_2484_ _2484_/A vssd1 vssd1 vccd1 vccd1 _4136_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4223_ _4222_/X _4415_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4223_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4154_ _4154_/A _4154_/B vssd1 vssd1 vccd1 vccd1 _4155_/B sky130_fd_sc_hd__or2_1
X_3105_ _3105_/A _3105_/B vssd1 vssd1 vccd1 vccd1 _3105_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4085_ _4085_/A vssd1 vssd1 vccd1 vccd1 _4085_/X sky130_fd_sc_hd__clkbuf_1
X_3036_ _3035_/X _2933_/A _2936_/B _2936_/D vssd1 vssd1 vccd1 vccd1 _3036_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2481__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3938_ _4451_/Q _3936_/X input3/X _3937_/X vssd1 vssd1 vccd1 vccd1 _4451_/D sky130_fd_sc_hd__a22o_1
X_3869_ _3869_/A vssd1 vssd1 vccd1 vccd1 _4488_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_39_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4347__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput28 addr_in[5] vssd1 vssd1 vccd1 vccd1 _2498_/A sky130_fd_sc_hd__buf_6
Xinput17 addr_in[24] vssd1 vssd1 vccd1 vccd1 _2537_/A sky130_fd_sc_hd__buf_6
Xinput39 data_in[15] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3426__S _3430_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3659__B1 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4257__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4772_ _4773_/CLK _4772_/D vssd1 vssd1 vccd1 vccd1 _4772_/Q sky130_fd_sc_hd__dfxtp_1
X_3723_ _4577_/Q _3717_/X _2493_/A _3718_/X vssd1 vssd1 vccd1 vccd1 _4577_/D sky130_fd_sc_hd__a22o_1
X_3654_ _3654_/A vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__clkbuf_2
X_2605_ _4624_/Q _2506_/X _4625_/Q _2508_/X vssd1 vssd1 vccd1 vccd1 _2605_/X sky130_fd_sc_hd__o22a_1
X_3585_ _3585_/A vssd1 vssd1 vccd1 vccd1 _4660_/D sky130_fd_sc_hd__clkbuf_1
X_2536_ _2536_/A vssd1 vssd1 vccd1 vccd1 _2536_/X sky130_fd_sc_hd__buf_2
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2467_ _2467_/A vssd1 vssd1 vccd1 vccd1 _4146_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4206_ _3977_/Y _3975_/A _4209_/S vssd1 vssd1 vccd1 vccd1 _4206_/X sky130_fd_sc_hd__mux2_1
X_2398_ _2390_/X _2391_/X _2393_/X _2397_/X vssd1 vssd1 vccd1 vccd1 _2403_/B sky130_fd_sc_hd__o211ai_1
XFILLER_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4137_ input7/X _4135_/Y _4145_/B vssd1 vssd1 vccd1 vccd1 _4137_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4068_ _4417_/X _4070_/B vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__and2_1
X_3019_ _2902_/A _3014_/X _2971_/B vssd1 vssd1 vccd1 vccd1 _3020_/B sky130_fd_sc_hd__a21bo_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3100__A _4571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__B1 _4387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output99_A _4513_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3370_ _3370_/A _4007_/B vssd1 vssd1 vccd1 vccd1 _3598_/C sky130_fd_sc_hd__nor2_1
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _4211_/X vssd1 vssd1 vccd1 vccd1 _2321_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3680__A _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _2471_/B _2418_/A _2413_/A _2413_/B vssd1 vssd1 vccd1 vccd1 _2355_/B sky130_fd_sc_hd__or4_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3280__A1 _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4755_ _4755_/CLK _4755_/D vssd1 vssd1 vccd1 vccd1 _4755_/Q sky130_fd_sc_hd__dfxtp_1
X_3706_ _4590_/Q _3703_/X input7/X _3704_/X vssd1 vssd1 vccd1 vccd1 _4590_/D sky130_fd_sc_hd__a22o_1
X_4686_ _4719_/CLK _4686_/D vssd1 vssd1 vccd1 vccd1 _4686_/Q sky130_fd_sc_hd__dfxtp_1
X_3637_ _4637_/Q _3633_/X _2455_/A _3634_/X vssd1 vssd1 vccd1 vccd1 _4637_/D sky130_fd_sc_hd__a22o_1
X_3568_ _4666_/Q _3559_/A _4262_/X _3560_/A vssd1 vssd1 vccd1 vccd1 _4666_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2519_ _2519_/A _2519_/B vssd1 vssd1 vccd1 vccd1 _2524_/C sky130_fd_sc_hd__nand2_1
X_3499_ _4698_/Q _3487_/A _4262_/X _3488_/A vssd1 vssd1 vccd1 vccd1 _4698_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4391__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3271__A1 _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3765__A _3772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4360__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3484__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input50_A data_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4382__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output137_A _3289_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3262__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2870_ input4/X _2971_/A _2851_/B _2869_/Y _2834_/X vssd1 vssd1 vccd1 vccd1 _2870_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4270__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4540_ _4769_/CLK _4540_/D vssd1 vssd1 vccd1 vccd1 _4540_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_10_clk clkbuf_opt_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4625_/CLK sky130_fd_sc_hd__clkbuf_16
X_4471_ _4531_/CLK _4471_/D vssd1 vssd1 vccd1 vccd1 _4471_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3422_ _4340_/X _4734_/Q _3586_/S vssd1 vssd1 vccd1 vccd1 _3423_/A sky130_fd_sc_hd__mux2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2525__B1 _2518_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3353_ _3974_/A _3972_/A _4020_/C _3581_/C vssd1 vssd1 vccd1 vccd1 _3572_/C sky130_fd_sc_hd__o211a_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2304_ _3104_/A _2290_/B _2301_/A _2301_/B vssd1 vssd1 vccd1 vccd1 _2305_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3284_ _3284_/A _3284_/B vssd1 vssd1 vccd1 vccd1 _3284_/X sky130_fd_sc_hd__and2_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4373__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2235_ _4585_/Q vssd1 vssd1 vccd1 vccd1 _2418_/A sky130_fd_sc_hd__inv_2
XFILLER_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3253__B2 _4547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3569__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2904__D _2949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4428__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2999_ _2998_/A _2998_/B _2998_/Y vssd1 vssd1 vccd1 vccd1 _3003_/A sky130_fd_sc_hd__a21oi_1
X_4738_ _4738_/CLK _4738_/D vssd1 vssd1 vccd1 vccd1 _4738_/Q sky130_fd_sc_hd__dfxtp_1
X_4669_ _4751_/CLK _4669_/D vssd1 vssd1 vccd1 vccd1 _4669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4355__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4419__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4103__B _4103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3434__S _3442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4265__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3971_ _3971_/A vssd1 vssd1 vccd1 vccd1 _3971_/Y sky130_fd_sc_hd__inv_2
X_2922_ _2923_/B vssd1 vssd1 vccd1 vccd1 _2922_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2853_ _4440_/Q vssd1 vssd1 vccd1 vccd1 _2853_/Y sky130_fd_sc_hd__inv_2
X_2784_ _2782_/C _2783_/Y _2776_/X vssd1 vssd1 vccd1 vccd1 _2785_/B sky130_fd_sc_hd__o21ai_1
X_4523_ _4771_/CLK _4523_/D vssd1 vssd1 vccd1 vccd1 _4523_/Q sky130_fd_sc_hd__dfxtp_2
X_4454_ _4589_/CLK _4454_/D vssd1 vssd1 vccd1 vccd1 _4454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4385_ _4625_/Q _4582_/Q _4547_/Q _4447_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4385_/X sky130_fd_sc_hd__mux4_2
X_3405_ _3405_/A vssd1 vssd1 vccd1 vccd1 _4743_/D sky130_fd_sc_hd__clkbuf_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ _4205_/X _3330_/Y _4354_/S _3335_/X vssd1 vssd1 vccd1 vccd1 _4761_/D sky130_fd_sc_hd__a31o_1
XFILLER_85_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3267_ _2803_/A _3098_/A _2543_/A _3105_/A vssd1 vssd1 vccd1 vccd1 _3276_/A sky130_fd_sc_hd__a22o_1
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ _4600_/Q vssd1 vssd1 vccd1 vccd1 _2273_/A sky130_fd_sc_hd__clkinv_2
X_3198_ _3198_/A _3198_/B vssd1 vssd1 vccd1 vccd1 _3198_/X sky130_fd_sc_hd__or2_1
XFILLER_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3299__B _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3701__A2 _3696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input13_A addr_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4414__A0 _4661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4170_ _4153_/A _4153_/B _4154_/B vssd1 vssd1 vccd1 vccd1 _4170_/X sky130_fd_sc_hd__a21bo_1
XFILLER_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3121_ _3121_/A _3121_/B vssd1 vssd1 vccd1 vccd1 _3121_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3052_ _4556_/Q vssd1 vssd1 vccd1 vccd1 _3116_/A sky130_fd_sc_hd__inv_2
XFILLER_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3954_ _4274_/X _4438_/Q _3960_/S vssd1 vssd1 vccd1 vccd1 _3955_/A sky130_fd_sc_hd__mux2_1
X_2905_ _2914_/B _2914_/D vssd1 vssd1 vccd1 vccd1 _2906_/B sky130_fd_sc_hd__or2_1
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3885_ _4223_/X _4480_/Q _3885_/S vssd1 vssd1 vccd1 vccd1 _3886_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2836_ _4449_/Q vssd1 vssd1 vccd1 vccd1 _3012_/A sky130_fd_sc_hd__inv_2
XANTENNA__4024__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2767_ _2737_/Y _2749_/X _2798_/A _2765_/A _2766_/Y vssd1 vssd1 vccd1 vccd1 _2767_/X
+ sky130_fd_sc_hd__o32a_1
X_2698_ _4639_/Q _2697_/Y _2694_/X vssd1 vssd1 vccd1 vccd1 _2698_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4506_ _4732_/CLK _4506_/D vssd1 vssd1 vccd1 vccd1 _4506_/Q sky130_fd_sc_hd__dfxtp_1
X_4437_ _4773_/CLK _4437_/D vssd1 vssd1 vccd1 vccd1 _4437_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input5_A addr_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4368_ _4755_/Q _4705_/Q _4672_/Q _4615_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4368_/X sky130_fd_sc_hd__mux4_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3319_/A vssd1 vssd1 vccd1 vccd1 _3320_/A sky130_fd_sc_hd__inv_2
X_4299_ _4104_/X _4431_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4299_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4411__A3 _4661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3670_ _3670_/A vssd1 vssd1 vccd1 vccd1 _4613_/D sky130_fd_sc_hd__clkbuf_1
X_2621_ _4646_/Q vssd1 vssd1 vccd1 vccd1 _2679_/A sky130_fd_sc_hd__inv_2
XANTENNA__3683__A _3697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput116 _4494_/Q vssd1 vssd1 vccd1 vccd1 data_out[21] sky130_fd_sc_hd__buf_2
X_2552_ _2549_/A _2551_/X _2549_/C vssd1 vssd1 vccd1 vccd1 _2552_/X sky130_fd_sc_hd__o21ba_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput105 _4484_/Q vssd1 vssd1 vccd1 vccd1 data_out[11] sky130_fd_sc_hd__buf_2
Xoutput138 _4695_/Q vssd1 vssd1 vccd1 vccd1 is_byte_out sky130_fd_sc_hd__buf_2
Xoutput127 _4504_/Q vssd1 vssd1 vccd1 vccd1 data_out[31] sky130_fd_sc_hd__buf_2
X_4222_ _4058_/X _4415_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4222_/X sky130_fd_sc_hd__mux2_1
X_2483_ input6/X vssd1 vssd1 vccd1 vccd1 _2484_/A sky130_fd_sc_hd__inv_2
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4153_ _4153_/A _4153_/B vssd1 vssd1 vccd1 vccd1 _4154_/B sky130_fd_sc_hd__or2_1
X_3104_ _3104_/A _3104_/B vssd1 vssd1 vccd1 vccd1 _3114_/A sky130_fd_sc_hd__nor2_1
X_4084_ _4423_/X _4092_/B vssd1 vssd1 vccd1 vccd1 _4085_/A sky130_fd_sc_hd__and2_1
X_3035_ _4347_/X _3035_/B vssd1 vssd1 vccd1 vccd1 _3035_/X sky130_fd_sc_hd__or2_1
XFILLER_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3937_ _3944_/A vssd1 vssd1 vccd1 vccd1 _3937_/X sky130_fd_sc_hd__clkbuf_2
X_3868_ _4326_/X _4488_/Q _3874_/S vssd1 vssd1 vccd1 vccd1 _3869_/A sky130_fd_sc_hd__mux2_1
X_2819_ _2819_/A _2884_/B _2819_/C _2819_/D vssd1 vssd1 vccd1 vccd1 _2819_/Y sky130_fd_sc_hd__nor4_1
X_3799_ _4526_/Q _3795_/X _4397_/X _3793_/X vssd1 vssd1 vccd1 vccd1 _4526_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4363__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 addr_in[25] vssd1 vssd1 vccd1 vccd1 _2816_/A sky130_fd_sc_hd__buf_8
Xinput29 addr_in[6] vssd1 vssd1 vccd1 vccd1 _2505_/A sky130_fd_sc_hd__buf_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2847__A _4447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3442__S _3442_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4273__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4771_ _4771_/CLK _4771_/D vssd1 vssd1 vccd1 vccd1 _4771_/Q sky130_fd_sc_hd__dfxtp_2
X_3722_ _4578_/Q _3717_/X _2492_/A _3718_/X vssd1 vssd1 vccd1 vccd1 _4578_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3653_ _4625_/Q _3647_/X _2507_/A _3648_/X vssd1 vssd1 vccd1 vccd1 _4625_/D sky130_fd_sc_hd__a22o_1
X_2604_ _2650_/A _2498_/A _2753_/A _2505_/A vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__o22a_1
X_3584_ _4213_/X _4660_/Q _3606_/S vssd1 vssd1 vccd1 vccd1 _3585_/A sky130_fd_sc_hd__mux2_1
X_2535_ _2535_/A vssd1 vssd1 vccd1 vccd1 _2536_/A sky130_fd_sc_hd__inv_2
X_2466_ _2466_/A vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4205_ _3963_/X _3290_/A _4354_/S vssd1 vssd1 vccd1 vccd1 _4205_/X sky130_fd_sc_hd__mux2_2
X_2397_ _3192_/A _2397_/B vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__or2_1
XFILLER_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _4136_/A _4136_/B _4136_/C vssd1 vssd1 vccd1 vccd1 _4145_/B sky130_fd_sc_hd__or3_2
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4067_ _4067_/A vssd1 vssd1 vccd1 vccd1 _4067_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3822__A1 _4509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3018_ _2412_/A _3013_/X _2409_/A _3017_/X vssd1 vssd1 vccd1 vccd1 _3026_/A sky130_fd_sc_hd__a22oi_1
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3822__B2 _3303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2492__A _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3588__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2561__B2 _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4358__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3510__A0 _4266_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3813__A1 _4516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _4357_/X _2315_/X _2317_/X _2319_/Y vssd1 vssd1 vccd1 vccd1 _2320_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2251_ _2251_/A _2399_/A vssd1 vssd1 vccd1 vccd1 _2413_/B sky130_fd_sc_hd__or2_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4268__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3900__S _3900_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_38_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3804__B2 _3800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3804__A1 _4523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4754_ _4755_/CLK _4754_/D vssd1 vssd1 vccd1 vccd1 _4754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _4591_/Q _3703_/X input8/X _3704_/X vssd1 vssd1 vccd1 vccd1 _4591_/D sky130_fd_sc_hd__a22o_1
X_4685_ _4740_/CLK _4685_/D vssd1 vssd1 vccd1 vccd1 _4685_/Q sky130_fd_sc_hd__dfxtp_1
X_3636_ _4638_/Q _3633_/X _2452_/A _3634_/X vssd1 vssd1 vccd1 vccd1 _4638_/D sky130_fd_sc_hd__a22o_1
X_3567_ _4667_/Q _3559_/A _4258_/X _3560_/A vssd1 vssd1 vccd1 vccd1 _4667_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3740__B1 _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2518_ _2478_/X _2489_/Y _2510_/X _2517_/X vssd1 vssd1 vccd1 vccd1 _2518_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__2487__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3498_ _4699_/Q _3487_/A _4258_/X _3488_/A vssd1 vssd1 vccd1 vccd1 _4699_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2449_ _2526_/A _4597_/Q _2824_/A _2256_/A vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__o22a_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4391__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4119_ _4119_/A _4119_/B vssd1 vssd1 vccd1 vccd1 _4120_/B sky130_fd_sc_hd__or2_1
XFILLER_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4220__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input43_A data_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4287__A1 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4382__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4470_ _4531_/CLK _4470_/D vssd1 vssd1 vccd1 vccd1 _4470_/Q sky130_fd_sc_hd__dfxtp_2
X_3421_ _3421_/A vssd1 vssd1 vccd1 vccd1 _4735_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3722__B1 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3352_ _3352_/A vssd1 vssd1 vccd1 vccd1 _3581_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2292_/X _2295_/Y _4346_/X _2296_/Y _2302_/Y vssd1 vssd1 vccd1 vccd1 _2305_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3283_ _3222_/X _3225_/Y _3282_/Y vssd1 vssd1 vccd1 vccd1 _3284_/B sky130_fd_sc_hd__o21bai_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4373__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2234_ _4586_/Q vssd1 vssd1 vccd1 vccd1 _2471_/B sky130_fd_sc_hd__inv_2
XFILLER_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4027__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2998_ _2998_/A _2998_/B vssd1 vssd1 vccd1 vccd1 _2998_/Y sky130_fd_sc_hd__nor2_1
X_4737_ _4737_/CLK _4737_/D vssd1 vssd1 vccd1 vccd1 _4737_/Q sky130_fd_sc_hd__dfxtp_1
X_4668_ _4750_/CLK _4668_/D vssd1 vssd1 vccd1 vccd1 _4668_/Q sky130_fd_sc_hd__dfxtp_1
X_3619_ _3655_/A vssd1 vssd1 vccd1 vccd1 _3634_/A sky130_fd_sc_hd__buf_4
X_4599_ _4600_/CLK _4599_/D vssd1 vssd1 vccd1 vccd1 _4599_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3713__B1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2516__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4269__A1 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3952__A0 _4266_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3180__A1 _4547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3970_ _3970_/A vssd1 vssd1 vccd1 vccd1 _3971_/A sky130_fd_sc_hd__clkbuf_2
X_2921_ _2921_/A _2926_/A _2926_/B vssd1 vssd1 vccd1 vccd1 _2923_/B sky130_fd_sc_hd__or3_1
XFILLER_62_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4281__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2852_ _4441_/Q vssd1 vssd1 vccd1 vccd1 _2852_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2783_ _2783_/A _2783_/B vssd1 vssd1 vccd1 vccd1 _2783_/Y sky130_fd_sc_hd__nor2_1
X_4522_ _4771_/CLK _4522_/D vssd1 vssd1 vccd1 vccd1 _4522_/Q sky130_fd_sc_hd__dfxtp_2
X_4453_ _4556_/CLK _4453_/D vssd1 vssd1 vccd1 vccd1 _4453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3404_ _4270_/X _4743_/Q _3408_/S vssd1 vssd1 vccd1 vccd1 _3405_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4384_ _4624_/Q _4581_/Q _4546_/Q _4446_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4384_/X sky130_fd_sc_hd__mux4_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3335_ _3329_/Y _4204_/X _3320_/X _2211_/A _4761_/Q vssd1 vssd1 vccd1 vccd1 _3335_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3266_ _2446_/A _4563_/Q _3228_/Y _3264_/X _3265_/X vssd1 vssd1 vccd1 vccd1 _3266_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2217_ _4601_/Q vssd1 vssd1 vccd1 vccd1 _2272_/B sky130_fd_sc_hd__clkinv_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _3196_/A _3196_/B _3198_/B vssd1 vssd1 vccd1 vccd1 _3197_/X sky130_fd_sc_hd__a21bo_1
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4191__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3934__B1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4111__B1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4366__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4414__A1 _4663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3925__B1 _2452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output74_A _4519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3120_ _4559_/Q _3118_/Y _3132_/B vssd1 vssd1 vccd1 vccd1 _3121_/B sky130_fd_sc_hd__o21ai_1
XFILLER_95_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3051_ _3051_/A _3137_/A _3130_/A vssd1 vssd1 vccd1 vccd1 _3132_/A sky130_fd_sc_hd__or3_1
XANTENNA__4276__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4405__A1 _4602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3953_ _3953_/A vssd1 vssd1 vccd1 vccd1 _4439_/D sky130_fd_sc_hd__clkbuf_1
X_2904_ _2904_/A _2939_/A _2938_/B _2949_/B vssd1 vssd1 vccd1 vccd1 _2914_/D sky130_fd_sc_hd__or4_2
XFILLER_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3884_ _3884_/A vssd1 vssd1 vccd1 vccd1 _4481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2835_ _4450_/Q vssd1 vssd1 vccd1 vccd1 _3014_/A sky130_fd_sc_hd__inv_2
X_2766_ _2761_/X _2762_/X _2765_/B _2765_/D vssd1 vssd1 vccd1 vccd1 _2766_/Y sky130_fd_sc_hd__a31oi_2
X_2697_ _2697_/A _2697_/B vssd1 vssd1 vccd1 vccd1 _2697_/Y sky130_fd_sc_hd__nor2_1
X_4505_ _4747_/CLK _4505_/D vssd1 vssd1 vccd1 vccd1 _4505_/Q sky130_fd_sc_hd__dfxtp_1
X_4436_ _4746_/CLK _4436_/D vssd1 vssd1 vccd1 vccd1 _4436_/Q sky130_fd_sc_hd__dfxtp_1
X_4367_ _4161_/X _2536_/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4367_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _3318_/A vssd1 vssd1 vccd1 vccd1 _3318_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4297_/X _4432_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__mux2_1
X_3249_ _2500_/A _3182_/A _2492_/A _3074_/A vssd1 vssd1 vccd1 vccd1 _3249_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4186__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4109__B _4109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4399__A0 _4639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ _4647_/Q vssd1 vssd1 vccd1 vccd1 _2674_/A sky130_fd_sc_hd__inv_2
XFILLER_9_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2551_ _2551_/A _2551_/B vssd1 vssd1 vccd1 vccd1 _2551_/X sky130_fd_sc_hd__and2_1
Xoutput106 _4485_/Q vssd1 vssd1 vccd1 vccd1 data_out[12] sky130_fd_sc_hd__buf_2
Xoutput128 _4476_/Q vssd1 vssd1 vccd1 vccd1 data_out[3] sky130_fd_sc_hd__buf_2
Xoutput139 _4185_/X vssd1 vssd1 vccd1 vccd1 is_data_to_cache sky130_fd_sc_hd__buf_2
X_2482_ _2482_/A vssd1 vssd1 vccd1 vccd1 _4136_/A sky130_fd_sc_hd__clkbuf_2
Xoutput117 _4495_/Q vssd1 vssd1 vccd1 vccd1 data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_5_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4221_ _4220_/X input34/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4221_/X sky130_fd_sc_hd__mux2_2
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4152_ _4152_/A _4152_/B vssd1 vssd1 vccd1 vccd1 _4153_/B sky130_fd_sc_hd__or2_1
XFILLER_68_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3103_ _4570_/Q _3099_/Y _4571_/Q _3100_/Y _3102_/X vssd1 vssd1 vccd1 vccd1 _3104_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4083_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4092_/B sky130_fd_sc_hd__buf_2
X_3034_ _2937_/A _2912_/X _2937_/C vssd1 vssd1 vccd1 vccd1 _3034_/X sky130_fd_sc_hd__o21ba_1
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3936_ _3943_/A vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3867_ _3867_/A vssd1 vssd1 vccd1 vccd1 _4489_/D sky130_fd_sc_hd__clkbuf_1
X_2818_ _2544_/A _4468_/Q _2546_/A _4467_/Q vssd1 vssd1 vccd1 vccd1 _2819_/D sky130_fd_sc_hd__a22o_1
X_3798_ _4527_/Q _3795_/X _4398_/X _3793_/X vssd1 vssd1 vccd1 vccd1 _4527_/D sky130_fd_sc_hd__a22o_1
X_2749_ _2744_/Y _2746_/X _2796_/D _2796_/C vssd1 vssd1 vccd1 vccd1 _2749_/X sky130_fd_sc_hd__o211a_1
X_4419_ _4734_/Q _4713_/Q _4680_/Q _4662_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4419_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 addr_in[26] vssd1 vssd1 vccd1 vccd1 _2815_/A sky130_fd_sc_hd__buf_6
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4400__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4770_ _4770_/CLK _4770_/D vssd1 vssd1 vccd1 vccd1 _4770_/Q sky130_fd_sc_hd__dfxtp_1
X_3721_ _4579_/Q _3717_/X _2500_/A _3718_/X vssd1 vssd1 vccd1 vccd1 _4579_/D sky130_fd_sc_hd__a22o_1
X_3652_ _4626_/Q _3647_/X _2472_/A _3648_/X vssd1 vssd1 vccd1 vccd1 _4626_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2603_ _4624_/Q vssd1 vssd1 vccd1 vccd1 _2753_/A sky130_fd_sc_hd__inv_2
X_3583_ _4367_/S _3328_/A _3582_/Y _4661_/Q _3582_/A vssd1 vssd1 vccd1 vccd1 _4661_/D
+ sky130_fd_sc_hd__a32o_1
X_2534_ _4158_/A _4604_/Q _4160_/A _4605_/Q vssd1 vssd1 vccd1 vccd1 _2550_/B sky130_fd_sc_hd__a22o_1
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2465_ _2465_/A vssd1 vssd1 vccd1 vccd1 _2466_/A sky130_fd_sc_hd__clkbuf_2
X_2396_ _2249_/A _2249_/B _2250_/B vssd1 vssd1 vccd1 vccd1 _2397_/B sky130_fd_sc_hd__a21bo_1
X_4204_ _3966_/X _4771_/Q _4354_/S vssd1 vssd1 vccd1 vccd1 _4204_/X sky130_fd_sc_hd__mux2_2
X_4135_ _4136_/B _4136_/C vssd1 vssd1 vccd1 vccd1 _4135_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ _4413_/X _4070_/B vssd1 vssd1 vccd1 vccd1 _4067_/A sky130_fd_sc_hd__and2_1
X_3017_ _2901_/A _2901_/B _3012_/B vssd1 vssd1 vccd1 vccd1 _3017_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__3822__A2 _3788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3588__B _4353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3919_ _4464_/Q _3915_/X _2537_/A _3916_/X vssd1 vssd1 vccd1 vccd1 _4464_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3274__B1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2250_ _2250_/A _2250_/B vssd1 vssd1 vccd1 vccd1 _2399_/A sky130_fd_sc_hd__or2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3689__A _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4284__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3804__A2 _3802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4753_ _4756_/CLK _4753_/D vssd1 vssd1 vccd1 vccd1 _4753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3704_ _3718_/A vssd1 vssd1 vccd1 vccd1 _3704_/X sky130_fd_sc_hd__clkbuf_2
X_4684_ _4747_/CLK _4684_/D vssd1 vssd1 vccd1 vccd1 _4684_/Q sky130_fd_sc_hd__dfxtp_1
X_3635_ _4639_/Q _3633_/X _2520_/A _3634_/X vssd1 vssd1 vccd1 vccd1 _4639_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4032__B _4032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3566_ _4668_/Q _3559_/A _4254_/X _3560_/A vssd1 vssd1 vccd1 vccd1 _4668_/D sky130_fd_sc_hd__a22o_1
X_3497_ _4367_/S _4354_/S _3496_/Y _4700_/Q _3496_/A vssd1 vssd1 vccd1 vccd1 _4700_/D
+ sky130_fd_sc_hd__a32o_1
X_2517_ input7/X _2255_/A _2485_/X _2516_/X vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__o22a_1
XFILLER_88_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2448_ _2448_/A vssd1 vssd1 vccd1 vccd1 _2526_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2379_ _2373_/Y _2377_/Y _4194_/X _2378_/B _2378_/Y vssd1 vssd1 vccd1 vccd1 _2379_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4118_ _4118_/A _4118_/B vssd1 vssd1 vccd1 vccd1 _4119_/B sky130_fd_sc_hd__or2_1
XFILLER_68_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4194__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4049_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4109_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input36_A data_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3798__A1 _4527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3420_ _4292_/X _4735_/Q _3420_/S vssd1 vssd1 vccd1 vccd1 _3421_/A sky130_fd_sc_hd__mux2_1
X_3351_ _3370_/A vssd1 vssd1 vccd1 vccd1 _3352_/A sky130_fd_sc_hd__inv_2
XANTENNA__4279__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2302_ _2302_/A vssd1 vssd1 vccd1 vccd1 _2302_/Y sky130_fd_sc_hd__inv_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _4762_/Q _3282_/B vssd1 vssd1 vccd1 vccd1 _3282_/Y sky130_fd_sc_hd__nand2_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2233_ _4587_/Q vssd1 vssd1 vccd1 vccd1 _2354_/A sky130_fd_sc_hd__inv_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3238__B1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3789__B2 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2997_ _3181_/A _2997_/B vssd1 vssd1 vccd1 vccd1 _3009_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4043__A _4375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4736_ _4736_/CLK _4736_/D vssd1 vssd1 vccd1 vccd1 _4736_/Q sky130_fd_sc_hd__dfxtp_1
X_4667_ _4706_/CLK _4667_/D vssd1 vssd1 vccd1 vccd1 _4667_/Q sky130_fd_sc_hd__dfxtp_1
X_3618_ _3654_/A vssd1 vssd1 vccd1 vccd1 _3655_/A sky130_fd_sc_hd__inv_4
XANTENNA__2498__A _2498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4598_ _4600_/CLK _4598_/D vssd1 vssd1 vccd1 vccd1 _4598_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3549_ _3549_/A vssd1 vssd1 vccd1 vccd1 _4677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_22_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_37_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4128__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2920_ _4468_/Q vssd1 vssd1 vccd1 vccd1 _2926_/A sky130_fd_sc_hd__inv_2
XFILLER_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2851_ _2851_/A _2851_/B _2851_/C _2851_/D vssd1 vssd1 vccd1 vccd1 _2851_/Y sky130_fd_sc_hd__nor4_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2782_ _2783_/B _2782_/B _2782_/C _2785_/A vssd1 vssd1 vccd1 vccd1 _2798_/C sky130_fd_sc_hd__or4_2
X_4521_ _4618_/CLK _4521_/D vssd1 vssd1 vccd1 vccd1 _4521_/Q sky130_fd_sc_hd__dfxtp_1
X_4452_ _4589_/CLK _4452_/D vssd1 vssd1 vccd1 vccd1 _4452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3403_ _3403_/A vssd1 vssd1 vccd1 vccd1 _4744_/D sky130_fd_sc_hd__clkbuf_1
X_4383_ _4623_/Q _4580_/Q _4545_/Q _4445_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4383_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ _3329_/Y _3330_/Y _4354_/S _3333_/X vssd1 vssd1 vccd1 vccd1 _4762_/D sky130_fd_sc_hd__a31o_1
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3265_ _2445_/A _4563_/Q _2526_/A _4562_/Q vssd1 vssd1 vccd1 vccd1 _3265_/X sky130_fd_sc_hd__a211o_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _4770_/Q vssd1 vssd1 vccd1 vccd1 _3290_/A sky130_fd_sc_hd__inv_2
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3196_ _3196_/A _3196_/B vssd1 vssd1 vccd1 vccd1 _3198_/B sky130_fd_sc_hd__or2_1
XFILLER_66_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3631__B1 _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4719_ _4719_/CLK _4719_/D vssd1 vssd1 vccd1 vccd1 _4719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3698__B1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4111__B2 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4111__A1 _3381_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2691__A _2702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4414__A2 _4665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3622__B1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3726__S _3780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3050_ _4560_/Q vssd1 vssd1 vccd1 vccd1 _3130_/A sky130_fd_sc_hd__inv_2
XFILLER_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3697__A _3697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4292__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3952_ _4266_/X _4439_/Q _3952_/S vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__mux2_1
X_2903_ _2967_/A _2967_/B _2903_/C _2971_/B vssd1 vssd1 vccd1 vccd1 _2949_/B sky130_fd_sc_hd__or4_4
X_3883_ _4219_/X _4481_/Q _3885_/S vssd1 vssd1 vccd1 vccd1 _3884_/A sky130_fd_sc_hd__mux2_1
X_2834_ input3/X _2902_/A vssd1 vssd1 vccd1 vccd1 _2834_/X sky130_fd_sc_hd__or2_1
X_2765_ _2765_/A _2765_/B _2765_/C _2765_/D vssd1 vssd1 vccd1 vccd1 _2798_/A sky130_fd_sc_hd__or4_4
X_4504_ _4752_/CLK _4504_/D vssd1 vssd1 vccd1 vccd1 _4504_/Q sky130_fd_sc_hd__dfxtp_1
X_2696_ _3134_/A _2706_/B _2340_/A _2695_/X vssd1 vssd1 vccd1 vccd1 _2709_/A sky130_fd_sc_hd__a22o_1
X_4435_ _4744_/CLK _4435_/D vssd1 vssd1 vccd1 vccd1 _4435_/Q sky130_fd_sc_hd__dfxtp_1
X_4366_ _4176_/X _4149_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4366_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _3314_/Y _3316_/A _3314_/A _3316_/Y _2212_/X vssd1 vssd1 vccd1 vccd1 _4766_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4106_/X _4432_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4297_/X sky130_fd_sc_hd__mux2_1
X_3248_ _3245_/X _3246_/X _3247_/X vssd1 vssd1 vccd1 vccd1 _3248_/X sky130_fd_sc_hd__a21bo_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3179_ _3179_/A _3179_/B vssd1 vssd1 vccd1 vccd1 _3179_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3852__A0 _4312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4399__A1 _4596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3310__A _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _2550_/A _2550_/B _2550_/C _2550_/D vssd1 vssd1 vccd1 vccd1 _2550_/X sky130_fd_sc_hd__or4_1
Xoutput107 _4486_/Q vssd1 vssd1 vccd1 vccd1 data_out[13] sky130_fd_sc_hd__buf_2
X_2481_ input7/X vssd1 vssd1 vccd1 vccd1 _2482_/A sky130_fd_sc_hd__inv_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput129 _4477_/Q vssd1 vssd1 vccd1 vccd1 data_out[4] sky130_fd_sc_hd__buf_2
Xoutput118 _4496_/Q vssd1 vssd1 vccd1 vccd1 data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4323__A1 _4372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4220_ _4013_/Y input34/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4220_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4151_ _4151_/A _4151_/B vssd1 vssd1 vccd1 vccd1 _4152_/B sky130_fd_sc_hd__or2_1
XANTENNA__4287__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3102_ _3102_/A _3102_/B vssd1 vssd1 vccd1 vccd1 _3102_/X sky130_fd_sc_hd__or2_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4082_ _4082_/A vssd1 vssd1 vccd1 vccd1 _4082_/X sky130_fd_sc_hd__clkbuf_1
X_3033_ _3033_/A vssd1 vssd1 vccd1 vccd1 _3033_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3935_ _4452_/Q _3929_/X input4/X _3930_/X vssd1 vssd1 vccd1 vccd1 _4452_/D sky130_fd_sc_hd__a22o_1
X_3866_ _4324_/X _4489_/Q _3874_/S vssd1 vssd1 vccd1 vccd1 _3867_/A sky130_fd_sc_hd__mux2_1
X_2817_ _4155_/A _4466_/Q _4154_/A _4465_/Q vssd1 vssd1 vccd1 vccd1 _2819_/C sky130_fd_sc_hd__a22o_1
X_3797_ _4528_/Q _3795_/X _4399_/X _3793_/X vssd1 vssd1 vccd1 vccd1 _4528_/D sky130_fd_sc_hd__a22o_1
X_2748_ _4187_/X _2748_/B vssd1 vssd1 vccd1 vccd1 _2796_/C sky130_fd_sc_hd__or2_1
X_2679_ _2679_/A _2679_/B vssd1 vssd1 vccd1 vccd1 _2679_/Y sky130_fd_sc_hd__nor2_1
X_4418_ _4733_/Q _4712_/Q _4679_/Q _4660_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4418_/X sky130_fd_sc_hd__mux4_1
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4349_ _4175_/A _4150_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4349_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input66_A is_byte vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2564__B1 _4637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4400__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2867__B2 _4447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3305__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3720_ _4580_/Q _3717_/X _2498_/A _3718_/X vssd1 vssd1 vccd1 vccd1 _4580_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_40_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4736_/CLK sky130_fd_sc_hd__clkbuf_16
X_3651_ _4627_/Q _3647_/X _2474_/A _3648_/X vssd1 vssd1 vccd1 vccd1 _4627_/D sky130_fd_sc_hd__a22o_1
X_2602_ _4623_/Q vssd1 vssd1 vccd1 vccd1 _2650_/A sky130_fd_sc_hd__inv_2
X_3582_ _3582_/A vssd1 vssd1 vccd1 vccd1 _3582_/Y sky130_fd_sc_hd__inv_2
X_2533_ _2533_/A vssd1 vssd1 vccd1 vccd1 _4160_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2464_ _2464_/A vssd1 vssd1 vccd1 vccd1 _2465_/A sky130_fd_sc_hd__inv_2
XFILLER_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2395_ _3008_/A vssd1 vssd1 vccd1 vccd1 _3192_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4203_ _3967_/Y _3962_/C _4338_/S vssd1 vssd1 vccd1 vccd1 _4203_/X sky130_fd_sc_hd__mux2_8
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4134_ _4134_/A _4134_/B vssd1 vssd1 vccd1 vccd1 _4136_/C sky130_fd_sc_hd__or2_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4065_ _4065_/A vssd1 vssd1 vccd1 vccd1 _4065_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3016_ _2412_/X _3013_/X _2417_/X _3015_/X vssd1 vssd1 vccd1 vccd1 _3026_/B sky130_fd_sc_hd__o22ai_1
XFILLER_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3918_ _4465_/Q _3915_/X _2816_/A _3916_/X vssd1 vssd1 vccd1 vccd1 _4465_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_31_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4740_/CLK sky130_fd_sc_hd__clkbuf_16
X_3849_ _3849_/A vssd1 vssd1 vccd1 vccd1 _4497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4394__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3274__A1 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4644_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4385__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4769_/CLK sky130_fd_sc_hd__clkbuf_16
X_4752_ _4752_/CLK _4752_/D vssd1 vssd1 vccd1 vccd1 _4752_/Q sky130_fd_sc_hd__dfxtp_1
X_3703_ _3717_/A vssd1 vssd1 vccd1 vccd1 _3703_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4683_ _4736_/CLK _4683_/D vssd1 vssd1 vccd1 vccd1 _4683_/Q sky130_fd_sc_hd__dfxtp_1
X_3634_ _3634_/A vssd1 vssd1 vccd1 vccd1 _3634_/X sky130_fd_sc_hd__clkbuf_2
X_3565_ _4669_/Q _3558_/X _4249_/X _3560_/X vssd1 vssd1 vccd1 vccd1 _4669_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3496_ _3496_/A vssd1 vssd1 vccd1 vccd1 _3496_/Y sky130_fd_sc_hd__inv_2
X_2516_ input6/X _2254_/A _2489_/A _2515_/X _2487_/X vssd1 vssd1 vccd1 vccd1 _2516_/X
+ sky130_fd_sc_hd__o221a_1
X_2447_ _2447_/A vssd1 vssd1 vccd1 vccd1 _2448_/A sky130_fd_sc_hd__inv_2
XANTENNA__4376__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2378_ _4194_/X _2378_/B vssd1 vssd1 vccd1 vccd1 _2378_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4117_ _4117_/A _4117_/B vssd1 vssd1 vccd1 vccd1 _4118_/B sky130_fd_sc_hd__or2_1
XFILLER_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_opt_2_0_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3256__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4048_ _4048_/A vssd1 vssd1 vccd1 vccd1 _4048_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input29_A addr_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3798__A2 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3350_ _3350_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _3370_/A sky130_fd_sc_hd__or2_1
X_2301_ _2301_/A _2301_/B vssd1 vssd1 vccd1 vccd1 _2302_/A sky130_fd_sc_hd__or2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3281_ _3266_/X _3276_/X _3280_/X vssd1 vssd1 vccd1 vccd1 _3282_/B sky130_fd_sc_hd__o21bai_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2232_ _4588_/Q vssd1 vssd1 vccd1 vccd1 _2487_/B sky130_fd_sc_hd__inv_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4752_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4295__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3238__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3789__A2 _3788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _4447_/Q _2995_/Y _2901_/B vssd1 vssd1 vccd1 vccd1 _2997_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4735_ _4735_/CLK _4735_/D vssd1 vssd1 vccd1 vccd1 _4735_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4043__B _4250_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4666_ _4706_/CLK _4666_/D vssd1 vssd1 vccd1 vccd1 _4666_/Q sky130_fd_sc_hd__dfxtp_1
X_3617_ _3633_/A vssd1 vssd1 vccd1 vccd1 _3617_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4597_ _4600_/CLK _4597_/D vssd1 vssd1 vccd1 vccd1 _4597_/Q sky130_fd_sc_hd__dfxtp_2
X_3548_ _4217_/X _4677_/Q _3548_/S vssd1 vssd1 vccd1 vccd1 _3549_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3479_ _3479_/A vssd1 vssd1 vccd1 vccd1 _4709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output135_A _4769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2850_ _2507_/A _2896_/A _2472_/A _2901_/A _2849_/X vssd1 vssd1 vccd1 vccd1 _2851_/D
+ sky130_fd_sc_hd__o221ai_1
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2781_ _2781_/A _2781_/B _2781_/C _2781_/D vssd1 vssd1 vccd1 vccd1 _2785_/A sky130_fd_sc_hd__or4_1
X_4520_ _4556_/CLK _4520_/D vssd1 vssd1 vccd1 vccd1 _4520_/Q sky130_fd_sc_hd__dfxtp_1
X_4451_ _4626_/CLK _4451_/D vssd1 vssd1 vccd1 vccd1 _4451_/Q sky130_fd_sc_hd__dfxtp_1
X_3402_ _4268_/X _4744_/Q _3408_/S vssd1 vssd1 vccd1 vccd1 _3403_/A sky130_fd_sc_hd__mux2_1
X_4382_ _4622_/Q _4579_/Q _4544_/Q _4444_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4382_/X sky130_fd_sc_hd__mux4_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _4205_/X _4204_/X _3320_/X _3962_/A _4762_/Q vssd1 vssd1 vccd1 vccd1 _3333_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_100_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3264_ _3263_/A _3233_/X _3259_/Y _3263_/X _3261_/X vssd1 vssd1 vccd1 vccd1 _3264_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _4772_/Q _4338_/S _2212_/X _3308_/A vssd1 vssd1 vccd1 vccd1 _4772_/D sky130_fd_sc_hd__o211a_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3163_/Y _3177_/X _3225_/A _3193_/A _3194_/Y vssd1 vssd1 vccd1 vccd1 _3195_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2979_ _2973_/X _2975_/X _3024_/B _3024_/D vssd1 vssd1 vccd1 vccd1 _2979_/Y sky130_fd_sc_hd__a31oi_1
X_4718_ _4740_/CLK _4718_/D vssd1 vssd1 vccd1 vccd1 _4718_/Q sky130_fd_sc_hd__dfxtp_1
X_4649_ _4649_/CLK _4649_/D vssd1 vssd1 vccd1 vccd1 _4649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3698__B2 _3697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3698__A1 _4596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4111__A2 _4013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3870__A1 _4487_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4414__A3 _4700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3386__A0 _4266_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4405__A3 _4467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3951_ _4440_/Q _3922_/A input1/X _3923_/A vssd1 vssd1 vccd1 vccd1 _4440_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2902_ _2902_/A _3014_/A _3012_/A _3012_/B vssd1 vssd1 vccd1 vccd1 _2971_/B sky130_fd_sc_hd__or4_2
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3882_ _3882_/A vssd1 vssd1 vccd1 vccd1 _4482_/D sky130_fd_sc_hd__clkbuf_1
X_2833_ _4451_/Q vssd1 vssd1 vccd1 vccd1 _2902_/A sky130_fd_sc_hd__inv_2
X_2764_ _2751_/A _2755_/B _3008_/A _2761_/B vssd1 vssd1 vccd1 vccd1 _2765_/D sky130_fd_sc_hd__a22o_1
X_4503_ _4732_/CLK _4503_/D vssd1 vssd1 vccd1 vccd1 _4503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2695_ _2645_/C _2694_/X _2692_/Y vssd1 vssd1 vccd1 vccd1 _2695_/X sky130_fd_sc_hd__a21o_1
X_4434_ _4730_/Q _4573_/Q _4611_/Q _4657_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4434_/X sky130_fd_sc_hd__mux4_1
X_4365_ _4144_/Y _2473_/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4365_/X sky130_fd_sc_hd__mux2_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _3316_/A vssd1 vssd1 vccd1 vccd1 _3316_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _4295_/X _4433_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4296_/X sky130_fd_sc_hd__mux2_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3247_ _4114_/A _4543_/Q _2494_/X _4542_/Q vssd1 vssd1 vccd1 vccd1 _3247_/X sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_21_clk_A clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4049__A _4094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3178_ _3178_/A _3182_/A _3182_/B vssd1 vssd1 vccd1 vccd1 _3179_/B sky130_fd_sc_hd__or3_1
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_36_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input11_A addr_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2207__A _3297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput119 _4497_/Q vssd1 vssd1 vccd1 vccd1 data_out[24] sky130_fd_sc_hd__buf_2
Xoutput108 _4487_/Q vssd1 vssd1 vccd1 vccd1 data_out[14] sky130_fd_sc_hd__buf_2
X_2480_ input3/X _2471_/B input2/X _2418_/A vssd1 vssd1 vccd1 vccd1 _2489_/B sky130_fd_sc_hd__a22o_1
XFILLER_49_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4150_ _4150_/A _4150_/B vssd1 vssd1 vccd1 vccd1 _4151_/B sky130_fd_sc_hd__or2_1
Xoutput90 _4534_/Q vssd1 vssd1 vccd1 vccd1 addr_out[27] sky130_fd_sc_hd__buf_2
X_3101_ _4570_/Q vssd1 vssd1 vccd1 vccd1 _3102_/A sky130_fd_sc_hd__inv_2
X_4081_ _4422_/X _4081_/B vssd1 vssd1 vccd1 vccd1 _4082_/A sky130_fd_sc_hd__and2_1
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3032_ _3032_/A _3032_/B _3032_/C _2963_/X vssd1 vssd1 vccd1 vccd1 _3041_/D sky130_fd_sc_hd__or4b_4
XFILLER_91_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3934_ _4453_/Q _3929_/X input5/X _3930_/X vssd1 vssd1 vccd1 vccd1 _4453_/D sky130_fd_sc_hd__a22o_1
X_3865_ _3887_/A vssd1 vssd1 vccd1 vccd1 _3874_/S sky130_fd_sc_hd__clkbuf_4
X_2816_ _2816_/A vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__inv_2
XFILLER_31_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3796_ _4529_/Q _3795_/X _4400_/X _3793_/X vssd1 vssd1 vccd1 vccd1 _4529_/D sky130_fd_sc_hd__a22o_1
X_2747_ _4192_/X _2747_/B vssd1 vssd1 vccd1 vccd1 _2796_/D sky130_fd_sc_hd__nand2_1
XANTENNA__4051__B _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2678_ _3104_/A _2678_/B vssd1 vssd1 vccd1 vccd1 _2689_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3770__B1 _2507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4417_ _4659_/Q _4711_/Q _4678_/Q _4613_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4417_/X sky130_fd_sc_hd__mux4_2
X_4348_ _4162_/Y _4160_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4348_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input3_A addr_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4279_ _4027_/Y input46/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4279_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3761__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2564__A1 _4638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input59_A data_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3305__B _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4241__A1 _3997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3650_ _4628_/Q _3647_/X input2/X _3648_/X vssd1 vssd1 vccd1 vccd1 _4628_/D sky130_fd_sc_hd__a22o_1
X_2601_ _2596_/X _2599_/X _2600_/X vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__a21bo_1
X_3581_ _4354_/X _4353_/X _3581_/C vssd1 vssd1 vccd1 vccd1 _3582_/A sky130_fd_sc_hd__or3_1
X_2532_ _2532_/A vssd1 vssd1 vccd1 vccd1 _2533_/A sky130_fd_sc_hd__inv_2
XANTENNA__3752__B1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4298__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3504__A0 _4264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4202_ _3968_/Y _3964_/Y _4338_/S vssd1 vssd1 vccd1 vccd1 _4202_/X sky130_fd_sc_hd__mux2_8
X_2463_ _4145_/A _4591_/Q _2467_/A _4592_/Q vssd1 vssd1 vccd1 vccd1 _2519_/B sky130_fd_sc_hd__o22a_1
XFILLER_87_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2394_ _4193_/X vssd1 vssd1 vccd1 vccd1 _3008_/A sky130_fd_sc_hd__inv_2
XFILLER_3_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4133_ _4133_/A _4133_/B vssd1 vssd1 vccd1 vccd1 _4134_/B sky130_fd_sc_hd__or2_1
X_4064_ _4412_/X _4070_/B vssd1 vssd1 vccd1 vccd1 _4065_/A sky130_fd_sc_hd__and2_1
X_3015_ _3014_/A _3014_/B _3014_/X vssd1 vssd1 vccd1 vccd1 _3015_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__2491__B1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4232__A1 _4005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3917_ _4466_/Q _3915_/X _2815_/A _3916_/X vssd1 vssd1 vccd1 vccd1 _4466_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3848_ _4308_/X _4497_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3849_/A sky130_fd_sc_hd__mux2_1
X_3779_ _4540_/Q _3750_/A input1/X _3751_/A vssd1 vssd1 vccd1 vccd1 _4540_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4394__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4385__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2220__A _4598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4214__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ _4751_/CLK _4751_/D vssd1 vssd1 vccd1 vccd1 _4751_/Q sky130_fd_sc_hd__dfxtp_1
X_4682_ _4736_/CLK _4682_/D vssd1 vssd1 vccd1 vccd1 _4682_/Q sky130_fd_sc_hd__dfxtp_1
X_3702_ _4592_/Q _3696_/X input9/X _3697_/X vssd1 vssd1 vccd1 vccd1 _4592_/D sky130_fd_sc_hd__a22o_1
X_3633_ _3633_/A vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3725__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3564_ _4670_/Q _3558_/X _4245_/X _3560_/X vssd1 vssd1 vccd1 vccd1 _4670_/D sky130_fd_sc_hd__a22o_1
X_3495_ _3569_/A _3576_/B _3581_/C vssd1 vssd1 vccd1 vccd1 _3496_/A sky130_fd_sc_hd__or3_1
X_2515_ input4/X _2355_/A _2489_/B _2514_/Y _2471_/X vssd1 vssd1 vccd1 vccd1 _2515_/X
+ sky130_fd_sc_hd__o221a_1
X_2446_ _2446_/A vssd1 vssd1 vccd1 vccd1 _4152_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4376__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2377_ _2377_/A vssd1 vssd1 vccd1 vccd1 _2377_/Y sky130_fd_sc_hd__inv_2
X_4116_ _3381_/D _4013_/A _2494_/X _4113_/Y vssd1 vssd1 vccd1 vccd1 _4116_/X sky130_fd_sc_hd__a31o_1
XFILLER_29_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4047_ _4377_/X _4250_/S vssd1 vssd1 vccd1 vccd1 _4048_/A sky130_fd_sc_hd__and2_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3716__B1 _2507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3835__S _3841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3707__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2300_ _4605_/Q _2285_/Y _2288_/X vssd1 vssd1 vccd1 vccd1 _2301_/B sky130_fd_sc_hd__o21ai_1
X_3280_ _2535_/A _3100_/Y _3269_/X _3279_/X vssd1 vssd1 vccd1 vccd1 _3280_/X sky130_fd_sc_hd__o22a_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _4589_/Q vssd1 vssd1 vccd1 vccd1 _2254_/A sky130_fd_sc_hd__inv_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3946__B1 _2498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2995_ _2995_/A _2995_/B vssd1 vssd1 vccd1 vccd1 _2995_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4734_ _4734_/CLK _4734_/D vssd1 vssd1 vccd1 vccd1 _4734_/Q sky130_fd_sc_hd__dfxtp_1
X_4665_ _4737_/CLK _4665_/D vssd1 vssd1 vccd1 vccd1 _4665_/Q sky130_fd_sc_hd__dfxtp_2
X_3616_ _3654_/A vssd1 vssd1 vccd1 vccd1 _3633_/A sky130_fd_sc_hd__clkbuf_4
X_4596_ _4639_/CLK _4596_/D vssd1 vssd1 vccd1 vccd1 _4596_/Q sky130_fd_sc_hd__dfxtp_2
X_3547_ _3547_/A vssd1 vssd1 vccd1 vccd1 _4678_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3478_ _4221_/X _4709_/Q _3482_/S vssd1 vssd1 vccd1 vccd1 _3479_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2429_ _2427_/C _2428_/X _2426_/X vssd1 vssd1 vccd1 vccd1 _2430_/B sky130_fd_sc_hd__o21ai_1
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input41_A data_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output128_A _4476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3928__B1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2780_ _2779_/X _2731_/X _2727_/X _2729_/X vssd1 vssd1 vccd1 vccd1 _2781_/C sky130_fd_sc_hd__o211ai_1
XFILLER_31_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _4626_/CLK _4450_/D vssd1 vssd1 vccd1 vccd1 _4450_/Q sky130_fd_sc_hd__dfxtp_1
X_4381_ _4621_/Q _4578_/Q _4543_/Q _4443_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4381_/X sky130_fd_sc_hd__mux4_1
X_3401_ _3401_/A vssd1 vssd1 vccd1 vccd1 _4745_/D sky130_fd_sc_hd__clkbuf_1
X_3332_ _4205_/X _4204_/X _4354_/S _3331_/X vssd1 vssd1 vccd1 vccd1 _4763_/D sky130_fd_sc_hd__a31o_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3263_/A _3263_/B _3263_/C _3263_/D vssd1 vssd1 vccd1 vccd1 _3263_/X sky130_fd_sc_hd__or4_1
X_3194_ _3192_/X _3186_/A _3188_/X _3193_/C vssd1 vssd1 vccd1 vccd1 _3194_/Y sky130_fd_sc_hd__a31oi_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _3962_/C _3965_/B vssd1 vssd1 vccd1 vccd1 _3308_/A sky130_fd_sc_hd__or2_1
XFILLER_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3919__B1 _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2978_ _2349_/A _2970_/B _2360_/X _2975_/B vssd1 vssd1 vccd1 vccd1 _3024_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4717_ _4738_/CLK _4717_/D vssd1 vssd1 vccd1 vccd1 _4717_/Q sky130_fd_sc_hd__dfxtp_1
X_4648_ _4649_/CLK _4648_/D vssd1 vssd1 vccd1 vccd1 _4648_/Q sky130_fd_sc_hd__dfxtp_2
X_4579_ _4623_/CLK _4579_/D vssd1 vssd1 vccd1 vccd1 _4579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3698__A2 _3696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4430__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3950_ _4441_/Q _3922_/A _3380_/A _3923_/A vssd1 vssd1 vccd1 vccd1 _4441_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2901_ _2901_/A _2901_/B vssd1 vssd1 vccd1 vccd1 _3012_/B sky130_fd_sc_hd__or2_1
X_3881_ _4338_/X _4482_/Q _3885_/S vssd1 vssd1 vccd1 vccd1 _3882_/A sky130_fd_sc_hd__mux2_1
X_2832_ _2967_/B vssd1 vssd1 vccd1 vccd1 _2971_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2763_ _2390_/X _2758_/X _2761_/X _2762_/X vssd1 vssd1 vccd1 vccd1 _2765_/C sky130_fd_sc_hd__o211ai_1
XFILLER_8_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4502_ _4629_/CLK _4502_/D vssd1 vssd1 vccd1 vccd1 _4502_/Q sky130_fd_sc_hd__dfxtp_2
X_2694_ _2694_/A _2697_/A _2697_/B vssd1 vssd1 vccd1 vccd1 _2694_/X sky130_fd_sc_hd__or3_1
X_4433_ _4731_/Q _4729_/Q _4697_/Q _4506_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4433_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4421__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4364_ _4143_/X _2513_/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4364_/X sky130_fd_sc_hd__mux2_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _4108_/X _4433_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4295_/X sky130_fd_sc_hd__mux2_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _2202_/C _3310_/B _4766_/Q _3325_/B vssd1 vssd1 vccd1 vccd1 _3316_/A sky130_fd_sc_hd__o22a_1
X_3246_ _2493_/A _3161_/A _3380_/A _3165_/Y vssd1 vssd1 vccd1 vccd1 _3246_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3234__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3172_/Y _3174_/X _3223_/D _3223_/C vssd1 vssd1 vccd1 vccd1 _3177_/X sky130_fd_sc_hd__o211a_1
XFILLER_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2812__B1 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4412__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2879__B1 _2873_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2983__A _4661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2207__B _2207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2223__A _4595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput109 _4488_/Q vssd1 vssd1 vccd1 vccd1 data_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__4403__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output72_A _4517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 _4535_/Q vssd1 vssd1 vccd1 vccd1 addr_out[28] sky130_fd_sc_hd__buf_2
XFILLER_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3100_ _4571_/Q vssd1 vssd1 vccd1 vccd1 _3100_/Y sky130_fd_sc_hd__inv_2
Xoutput80 _4525_/Q vssd1 vssd1 vccd1 vccd1 addr_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__3989__A _3989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4080_ _4080_/A vssd1 vssd1 vccd1 vccd1 _4080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3031_ _3031_/A _3031_/B vssd1 vssd1 vccd1 vccd1 _3032_/B sky130_fd_sc_hd__or2_1
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3933_ _4454_/Q _3929_/X input6/X _3930_/X vssd1 vssd1 vccd1 vccd1 _4454_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3864_ _3864_/A vssd1 vssd1 vccd1 vccd1 _4490_/D sky130_fd_sc_hd__clkbuf_1
X_2815_ _2815_/A vssd1 vssd1 vccd1 vccd1 _4155_/A sky130_fd_sc_hd__clkinv_4
XFILLER_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3795_ _3816_/A vssd1 vssd1 vccd1 vccd1 _3795_/X sky130_fd_sc_hd__buf_4
X_2746_ _4187_/X _2748_/B vssd1 vssd1 vccd1 vccd1 _2746_/X sky130_fd_sc_hd__and2_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2677_ _4648_/Q _2675_/Y _4649_/Q _2625_/Y _2676_/X vssd1 vssd1 vccd1 vccd1 _2678_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3770__A1 _4547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4416_ _4374_/X _4373_/X _4372_/X _4369_/X input1/X _3380_/A vssd1 vssd1 vccd1 vccd1
+ _4416_/X sky130_fd_sc_hd__mux4_1
X_4347_ _4183_/A _2803_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4347_/X sky130_fd_sc_hd__mux2_2
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4278_ _4277_/X input47/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4278_/X sky130_fd_sc_hd__mux2_1
X_3229_ _2454_/A _4560_/Q _2457_/A _4559_/Q vssd1 vssd1 vccd1 vccd1 _3263_/A sky130_fd_sc_hd__a22o_1
XFILLER_100_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3038__B1 _3029_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2600_ _4623_/Q _2499_/X _4622_/Q _2501_/X vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__o22a_1
XFILLER_61_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3580_ _3580_/A vssd1 vssd1 vccd1 vccd1 _4662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2531_ _2531_/A vssd1 vssd1 vccd1 vccd1 _4158_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_35_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4201_ _3982_/Y _3981_/A _4209_/S vssd1 vssd1 vccd1 vccd1 _4201_/X sky130_fd_sc_hd__mux2_1
X_2462_ _2462_/A vssd1 vssd1 vccd1 vccd1 _2467_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2393_ _2762_/A _2393_/B vssd1 vssd1 vccd1 vccd1 _2393_/X sky130_fd_sc_hd__or2_1
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4132_ _4132_/A _4132_/B vssd1 vssd1 vccd1 vccd1 _4133_/B sky130_fd_sc_hd__or2_1
XFILLER_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _4063_/A vssd1 vssd1 vccd1 vccd1 _4063_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3014_ _3014_/A _3014_/B vssd1 vssd1 vccd1 vccd1 _3014_/X sky130_fd_sc_hd__or2_1
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2491__A1 _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3916_ _3923_/A vssd1 vssd1 vccd1 vccd1 _3916_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4062__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3847_ _3847_/A vssd1 vssd1 vccd1 vccd1 _4498_/D sky130_fd_sc_hd__clkbuf_1
X_3778_ _4541_/Q _3750_/A _3380_/A _3751_/A vssd1 vssd1 vccd1 vccd1 _4541_/D sky130_fd_sc_hd__a22o_1
XANTENNA__2798__A _2798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2729_ _3156_/A _2729_/B vssd1 vssd1 vccd1 vccd1 _2729_/X sky130_fd_sc_hd__or2_1
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4750_ _4750_/CLK _4750_/D vssd1 vssd1 vccd1 vccd1 _4750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4681_ _4733_/CLK _4681_/D vssd1 vssd1 vccd1 vccd1 _4681_/Q sky130_fd_sc_hd__dfxtp_1
X_3701_ _4593_/Q _3696_/X _2464_/A _3697_/X vssd1 vssd1 vccd1 vccd1 _4593_/D sky130_fd_sc_hd__a22o_1
X_3632_ _4640_/Q _3626_/X _2447_/A _3627_/X vssd1 vssd1 vccd1 vccd1 _4640_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3725__B2 _3697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2528__A2 _4598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3563_ _4671_/Q _3558_/X _4241_/X _3560_/X vssd1 vssd1 vccd1 vccd1 _4671_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3494_ _4701_/Q _3487_/A _4254_/X _3488_/A vssd1 vssd1 vccd1 vccd1 _4701_/D sky130_fd_sc_hd__a22o_1
X_2514_ _2512_/X _4585_/Q _2513_/X _4584_/Q _2476_/X vssd1 vssd1 vccd1 vccd1 _2514_/Y
+ sky130_fd_sc_hd__a221oi_2
XFILLER_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2445_ _2445_/A vssd1 vssd1 vccd1 vccd1 _2446_/A sky130_fd_sc_hd__clkbuf_2
X_4115_ _2492_/A _4113_/Y _4117_/B vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__o21a_1
X_2376_ input1/X _4367_/S _4014_/A _3381_/B vssd1 vssd1 vccd1 vccd1 _2377_/A sky130_fd_sc_hd__o22a_4
XANTENNA__3242__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4057__B _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4046_ _4046_/A vssd1 vssd1 vccd1 vccd1 _4046_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3661__B1 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3652__B1 _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _4590_/Q vssd1 vssd1 vccd1 vccd1 _2255_/A sky130_fd_sc_hd__inv_2
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3997__A _3997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3643__B1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2994_ _2994_/A _2998_/A _2998_/B vssd1 vssd1 vccd1 vccd1 _2995_/B sky130_fd_sc_hd__or3_1
XANTENNA__4199__A1 _3989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4733_ _4733_/CLK _4733_/D vssd1 vssd1 vccd1 vccd1 _4733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4664_ _4733_/CLK _4664_/D vssd1 vssd1 vccd1 vccd1 _4664_/Q sky130_fd_sc_hd__dfxtp_1
X_4595_ _4639_/CLK _4595_/D vssd1 vssd1 vccd1 vccd1 _4595_/Q sky130_fd_sc_hd__dfxtp_2
X_3615_ _3965_/A _3615_/B vssd1 vssd1 vccd1 vccd1 _3654_/A sky130_fd_sc_hd__or2_4
X_3546_ _4215_/X _4678_/Q _3548_/S vssd1 vssd1 vccd1 vccd1 _3547_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3477_ _3477_/A vssd1 vssd1 vccd1 vccd1 _4710_/D sky130_fd_sc_hd__clkbuf_1
X_2428_ _2415_/Y _2428_/B vssd1 vssd1 vccd1 vccd1 _2428_/X sky130_fd_sc_hd__and2b_1
XFILLER_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2359_ _4355_/X vssd1 vssd1 vccd1 vccd1 _3156_/A sky130_fd_sc_hd__inv_2
XFILLER_28_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4029_ input1/X _4039_/B _4029_/C vssd1 vssd1 vccd1 vccd1 _4029_/Y sky130_fd_sc_hd__nor3_1
XFILLER_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3846__S _3852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_A data_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3625__B1 _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4380_ _4620_/Q _4577_/Q _4542_/Q _4442_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4380_/X sky130_fd_sc_hd__mux4_1
X_3400_ _4280_/X _4745_/Q _3412_/S vssd1 vssd1 vccd1 vccd1 _3401_/A sky130_fd_sc_hd__mux2_1
X_3331_ _3329_/Y _3330_/Y _3320_/X _3962_/A _4763_/Q vssd1 vssd1 vccd1 vccd1 _3331_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_98_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ input8/X _3116_/A _3261_/X vssd1 vssd1 vccd1 vccd1 _3263_/D sky130_fd_sc_hd__o21ai_1
XFILLER_100_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3193_ _3193_/A _3193_/B _3193_/C _3192_/X vssd1 vssd1 vccd1 vccd1 _3225_/A sky130_fd_sc_hd__or4b_2
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _4772_/Q vssd1 vssd1 vccd1 vccd1 _3962_/C sky130_fd_sc_hd__clkinv_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3520__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2977_ _2353_/X _2973_/B _2779_/X _2976_/X vssd1 vssd1 vccd1 vccd1 _3024_/B sky130_fd_sc_hd__a22o_1
X_4716_ _4737_/CLK _4716_/D vssd1 vssd1 vccd1 vccd1 _4716_/Q sky130_fd_sc_hd__dfxtp_1
X_4647_ _4649_/CLK _4647_/D vssd1 vssd1 vccd1 vccd1 _4647_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4070__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4578_ _4621_/CLK _4578_/D vssd1 vssd1 vccd1 vccd1 _4578_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3529_ _3529_/A vssd1 vssd1 vccd1 vccd1 _4686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4430__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output140_A _3341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2900_ _2994_/A _2998_/A _2900_/C _2998_/B vssd1 vssd1 vccd1 vccd1 _2901_/B sky130_fd_sc_hd__or4_2
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3880_ _3880_/A vssd1 vssd1 vccd1 vccd1 _4483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2831_ _4452_/Q vssd1 vssd1 vccd1 vccd1 _2967_/B sky130_fd_sc_hd__inv_2
XFILLER_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2762_ _2762_/A _2762_/B vssd1 vssd1 vccd1 vccd1 _2762_/X sky130_fd_sc_hd__or2_1
XFILLER_8_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4501_ _4693_/CLK _4501_/D vssd1 vssd1 vccd1 vccd1 _4501_/Q sky130_fd_sc_hd__dfxtp_4
X_2693_ _4641_/Q _2692_/Y _2668_/D vssd1 vssd1 vccd1 vccd1 _2706_/B sky130_fd_sc_hd__o21ai_1
X_4432_ _4732_/Q _4728_/Q _4696_/Q _4658_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4432_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4421__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4363_ _4177_/X _4148_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4363_/X sky130_fd_sc_hd__mux2_2
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _4293_/X _4434_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4294_/X sky130_fd_sc_hd__mux2_1
X_3314_ _3314_/A vssd1 vssd1 vccd1 vccd1 _3314_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3245_ _3380_/A _3165_/Y input1/X _3164_/Y vssd1 vssd1 vccd1 vccd1 _3245_/X sky130_fd_sc_hd__a211o_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3176_ _4187_/X _3176_/B vssd1 vssd1 vccd1 vccd1 _3223_/C sky130_fd_sc_hd__or2_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2812__A1 _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4412__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4403__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 _4536_/Q vssd1 vssd1 vccd1 vccd1 addr_out[29] sky130_fd_sc_hd__buf_2
XFILLER_68_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput81 _4526_/Q vssd1 vssd1 vccd1 vccd1 addr_out[19] sky130_fd_sc_hd__buf_2
X_3030_ _2317_/X _2961_/X _2962_/Y vssd1 vssd1 vccd1 vccd1 _3031_/B sky130_fd_sc_hd__o21ai_1
XFILLER_63_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3932_ _4455_/Q _3929_/X input7/X _3930_/X vssd1 vssd1 vccd1 vccd1 _4455_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_43_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4770_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_9_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3863_ _4322_/X _4490_/Q _3863_/S vssd1 vssd1 vccd1 vccd1 _3864_/A sky130_fd_sc_hd__mux2_1
X_2814_ _2537_/A _2914_/B _2816_/A _2914_/A vssd1 vssd1 vccd1 vccd1 _2884_/B sky130_fd_sc_hd__a22o_1
X_3794_ _4530_/Q _3788_/X _4401_/X _3793_/X vssd1 vssd1 vccd1 vccd1 _4530_/D sky130_fd_sc_hd__a22o_1
X_2745_ _2735_/A _2735_/B _2735_/Y vssd1 vssd1 vccd1 vccd1 _2748_/B sky130_fd_sc_hd__a21oi_1
X_2676_ _2676_/A _2676_/B vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__or2_1
X_4415_ _4756_/Q _4706_/Q _4673_/Q _4608_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4415_/X sky130_fd_sc_hd__mux4_2
X_4346_ _4164_/X _4157_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4346_/X sky130_fd_sc_hd__mux2_4
XFILLER_100_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4277_ _4028_/Y input47/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4277_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3228_ _2520_/A _3137_/A _3227_/X vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3159_ _2349_/A _3150_/B _2360_/X _3156_/B vssd1 vssd1 vccd1 vccd1 _3208_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3038__B2 _3041_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2308__B _2318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4733_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4397__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4639_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2530_ _2803_/A vssd1 vssd1 vccd1 vccd1 _2531_/A sky130_fd_sc_hd__inv_2
XANTENNA__4388__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2461_ input9/X vssd1 vssd1 vccd1 vccd1 _2462_/A sky130_fd_sc_hd__inv_2
X_4200_ _3986_/Y _3985_/A _4209_/S vssd1 vssd1 vccd1 vccd1 _4200_/X sky130_fd_sc_hd__mux2_1
X_2392_ _2762_/A _2393_/B _2390_/X _2391_/X vssd1 vssd1 vccd1 vccd1 _2403_/A sky130_fd_sc_hd__a22o_1
X_4131_ _4131_/A _4131_/B vssd1 vssd1 vccd1 vccd1 _4132_/B sky130_fd_sc_hd__or2_1
XFILLER_95_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4062_ _4371_/X _4070_/B vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__and2_1
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3013_ _3012_/A _3012_/B _3014_/B vssd1 vssd1 vccd1 vccd1 _3013_/X sky130_fd_sc_hd__a21bo_1
XFILLER_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_16_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4618_/CLK sky130_fd_sc_hd__clkbuf_16
X_3915_ _3922_/A vssd1 vssd1 vccd1 vccd1 _3915_/X sky130_fd_sc_hd__clkbuf_2
X_3846_ _4306_/X _4498_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__mux2_1
X_3777_ _4542_/Q _3771_/X _2493_/A _3772_/X vssd1 vssd1 vccd1 vccd1 _4542_/D sky130_fd_sc_hd__a22o_1
X_2728_ _2722_/A _2722_/B _2722_/Y vssd1 vssd1 vccd1 vccd1 _2729_/B sky130_fd_sc_hd__a21o_1
XANTENNA__4379__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2659_ _2668_/B _2668_/D vssd1 vssd1 vccd1 vccd1 _2660_/B sky130_fd_sc_hd__or2_1
XFILLER_101_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4329_ _4071_/X _4418_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4329_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3703__A _3717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3584__S _3606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A data_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3700_ _4594_/Q _3696_/X _2455_/A _3697_/X vssd1 vssd1 vccd1 vccd1 _4594_/D sky130_fd_sc_hd__a22o_1
X_4680_ _4719_/CLK _4680_/D vssd1 vssd1 vccd1 vccd1 _4680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3631_ _4641_/Q _3626_/X _2824_/A _3627_/X vssd1 vssd1 vccd1 vccd1 _4641_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3725__A2 _3696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3562_ _4672_/Q _3558_/X _4237_/X _3560_/X vssd1 vssd1 vccd1 vccd1 _4672_/D sky130_fd_sc_hd__a22o_1
X_2513_ _2513_/A vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__clkbuf_2
X_3493_ _4702_/Q _3486_/X _4249_/X _3488_/X vssd1 vssd1 vccd1 vccd1 _4702_/D sky130_fd_sc_hd__a22o_1
X_2444_ _2824_/A vssd1 vssd1 vccd1 vccd1 _2445_/A sky130_fd_sc_hd__clkinv_2
Xclkbuf_leaf_5_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4773_/CLK sky130_fd_sc_hd__clkbuf_16
X_2375_ _4367_/S vssd1 vssd1 vccd1 vccd1 _3381_/B sky130_fd_sc_hd__inv_2
XFILLER_96_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4114_ _4114_/A _4114_/B vssd1 vssd1 vccd1 vccd1 _4117_/B sky130_fd_sc_hd__or2_1
XFILLER_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4045_ _4376_/X _4250_/S vssd1 vssd1 vccd1 vccd1 _4046_/A sky130_fd_sc_hd__and2_1
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3661__B2 _3634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4073__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2767__A3 _2798_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3829_ _2204_/Y _3342_/B _4195_/S vssd1 vssd1 vccd1 vccd1 _3830_/B sky130_fd_sc_hd__o21a_1
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3652__B2 _3648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3579__S _3606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_34_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_49_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4203__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3343__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2993_ _2988_/X _3039_/B _2991_/Y _2992_/X vssd1 vssd1 vccd1 vccd1 _2993_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4732_ _4732_/CLK _4732_/D vssd1 vssd1 vccd1 vccd1 _4732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4663_ _4737_/CLK _4663_/D vssd1 vssd1 vccd1 vccd1 _4663_/Q sky130_fd_sc_hd__dfxtp_4
X_3614_ _3614_/A vssd1 vssd1 vccd1 vccd1 _4650_/D sky130_fd_sc_hd__clkbuf_1
X_4594_ _4637_/CLK _4594_/D vssd1 vssd1 vccd1 vccd1 _4594_/Q sky130_fd_sc_hd__dfxtp_2
X_3545_ _3545_/A vssd1 vssd1 vccd1 vccd1 _4679_/D sky130_fd_sc_hd__clkbuf_1
X_3476_ _4217_/X _4710_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3477_/A sky130_fd_sc_hd__mux2_1
X_2427_ _2430_/A _2427_/B _2427_/C _2426_/X vssd1 vssd1 vccd1 vccd1 _2443_/C sky130_fd_sc_hd__or4b_2
XFILLER_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2358_ _2353_/X _2356_/Y _4359_/X _2357_/Y vssd1 vssd1 vccd1 vccd1 _2358_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4068__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2289_ _4605_/Q _2285_/Y _4606_/Q _2286_/Y _2288_/X vssd1 vssd1 vccd1 vccd1 _2290_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4028_ input1/X _4038_/B _4029_/C vssd1 vssd1 vccd1 vccd1 _4028_/Y sky130_fd_sc_hd__nor3_1
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input27_A addr_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2507__A _2507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output95_A _4538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3330_ _4204_/X vssd1 vssd1 vccd1 vccd1 _3330_/Y sky130_fd_sc_hd__inv_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _2521_/A _4561_/Q _2453_/A _4560_/Q vssd1 vssd1 vccd1 vccd1 _3261_/X sky130_fd_sc_hd__o22a_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3192_ _3192_/A _3192_/B vssd1 vssd1 vccd1 vccd1 _3192_/X sky130_fd_sc_hd__or2_1
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _3962_/A vssd1 vssd1 vccd1 vccd1 _2212_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4408__A3 _4470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3520__B _3556_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2976_ _2971_/A _2971_/B _2971_/Y vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__a21o_1
X_4715_ _4736_/CLK _4715_/D vssd1 vssd1 vccd1 vccd1 _4715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4646_ _4649_/CLK _4646_/D vssd1 vssd1 vccd1 vccd1 _4646_/Q sky130_fd_sc_hd__dfxtp_2
X_4577_ _4621_/CLK _4577_/D vssd1 vssd1 vccd1 vccd1 _4577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3528_ _4282_/X _4686_/Q _3530_/S vssd1 vssd1 vccd1 vccd1 _3529_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3459_ _3459_/A vssd1 vssd1 vccd1 vccd1 _4718_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3304__B1 _3303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3855__A1 _4494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3711__A _3718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4280__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3857__S _3863_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2594__B2 _3380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3846__A1 _4498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4271__A1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2830_ _2874_/B _2878_/B _2874_/A vssd1 vssd1 vccd1 vccd1 _2830_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2761_ _3008_/A _2761_/B vssd1 vssd1 vccd1 vccd1 _2761_/X sky130_fd_sc_hd__or2_1
XFILLER_12_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2692_ _2692_/A _2697_/B vssd1 vssd1 vccd1 vccd1 _2692_/Y sky130_fd_sc_hd__nor2_1
X_4500_ _4693_/CLK _4500_/D vssd1 vssd1 vccd1 vccd1 _4500_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4431_ _4752_/Q _4727_/Q _4694_/Q _4439_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4431_/X sky130_fd_sc_hd__mux4_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4362_ _4172_/X _4151_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4362_/X sky130_fd_sc_hd__mux2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _4110_/X _4434_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4293_/X sky130_fd_sc_hd__mux2_1
X_3313_ _2202_/A _3310_/B _3319_/A _3318_/A vssd1 vssd1 vccd1 vccd1 _3314_/A sky130_fd_sc_hd__o211a_1
X_3244_ _3244_/A _3244_/B _3244_/C _3244_/D vssd1 vssd1 vccd1 vccd1 _3244_/Y sky130_fd_sc_hd__nor4_1
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3837__A1 _4502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3175_ _4192_/X _3175_/B vssd1 vssd1 vccd1 vccd1 _3223_/D sky130_fd_sc_hd__nand2_1
XFILLER_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2959_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2959_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4081__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3773__B1 _2505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2576__B2 _2474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4629_ _4629_/CLK _4629_/D vssd1 vssd1 vccd1 vccd1 _4629_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4301__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4253__A1 _3985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2567__A1 _4637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3616__A _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2520__A _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4211__S _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput93 _4509_/Q vssd1 vssd1 vccd1 vccd1 addr_out[2] sky130_fd_sc_hd__buf_2
Xoutput82 _4508_/Q vssd1 vssd1 vccd1 vccd1 addr_out[1] sky130_fd_sc_hd__buf_2
Xoutput71 _4507_/Q vssd1 vssd1 vccd1 vccd1 addr_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__3819__A1 _4512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3819__B2 _3814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4244__A1 _3993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3931_ _4456_/Q _3929_/X input8/X _3930_/X vssd1 vssd1 vccd1 vccd1 _4456_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3862_ _3862_/A vssd1 vssd1 vccd1 vccd1 _4491_/D sky130_fd_sc_hd__clkbuf_1
X_2813_ _4465_/Q vssd1 vssd1 vccd1 vccd1 _2914_/A sky130_fd_sc_hd__inv_2
X_3793_ _3814_/A vssd1 vssd1 vccd1 vccd1 _3793_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3755__B1 _2464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2744_ _4194_/X _2742_/B _2743_/X vssd1 vssd1 vccd1 vccd1 _2744_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2675_ _2676_/B vssd1 vssd1 vccd1 vccd1 _2675_/Y sky130_fd_sc_hd__inv_2
X_4414_ _4661_/Q _4663_/Q _4665_/Q _4700_/Q _4042_/Y _3971_/A vssd1 vssd1 vccd1 vccd1
+ _4414_/X sky130_fd_sc_hd__mux4_2
X_4345_ _4170_/X _4153_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4345_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4276_ _4275_/X input48/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4276_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3227_ _2445_/A _4563_/Q _2447_/A _3051_/A _3226_/X vssd1 vssd1 vccd1 vccd1 _3227_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3158_ _2353_/X _3154_/B _2779_/X _3157_/X vssd1 vssd1 vccd1 vccd1 _3208_/B sky130_fd_sc_hd__a22o_1
XFILLER_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _3089_/A _3089_/B vssd1 vssd1 vccd1 vccd1 _3090_/C sky130_fd_sc_hd__or2_1
XFILLER_23_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2797__A1 _2377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3746__B1 _2816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4397__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3870__S _3874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2485__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4388__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3346__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2460_ _2460_/A vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__clkbuf_2
X_2391_ _2247_/A _2247_/B _2248_/B vssd1 vssd1 vccd1 vccd1 _2391_/X sky130_fd_sc_hd__a21bo_1
X_4130_ _4130_/A _4130_/B vssd1 vssd1 vccd1 vccd1 _4131_/B sky130_fd_sc_hd__or2_1
XANTENNA__3780__S _3780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4061_ _4109_/B vssd1 vssd1 vccd1 vccd1 _4070_/B sky130_fd_sc_hd__buf_2
XFILLER_1_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3012_ _3012_/A _3012_/B vssd1 vssd1 vccd1 vccd1 _3014_/B sky130_fd_sc_hd__or2_1
XFILLER_36_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4217__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3914_ _4467_/Q _3906_/X _2545_/A _3909_/X vssd1 vssd1 vccd1 vccd1 _4467_/D sky130_fd_sc_hd__a22o_1
XANTENNA__3728__A0 _4256_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3845_ _3845_/A vssd1 vssd1 vccd1 vccd1 _4499_/D sky130_fd_sc_hd__clkbuf_1
X_3776_ _4543_/Q _3771_/X _2492_/A _3772_/X vssd1 vssd1 vccd1 vccd1 _4543_/D sky130_fd_sc_hd__a22o_1
X_2727_ _3154_/A _2727_/B vssd1 vssd1 vccd1 vccd1 _2727_/X sky130_fd_sc_hd__or2_1
XANTENNA__2798__C _2798_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4379__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2658_ _2658_/A _2692_/A _2691_/B _2702_/B vssd1 vssd1 vccd1 vccd1 _2668_/D sky130_fd_sc_hd__or4_2
X_2589_ _2589_/A _2589_/B _2589_/C _2589_/D vssd1 vssd1 vccd1 vccd1 _2589_/Y sky130_fd_sc_hd__nor4_1
X_4328_ _4327_/X _4419_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4328_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input1_A addr_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4259_ _4038_/Y input56/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4259_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3719__B1 _2505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3166__A _4663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input57_A data_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_0_0_clk_A clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3630_ _4642_/Q _3626_/X _2537_/A _3627_/X vssd1 vssd1 vccd1 vccd1 _4642_/D sky130_fd_sc_hd__a22o_1
X_3561_ _4673_/Q _3558_/X _4233_/X _3560_/X vssd1 vssd1 vccd1 vccd1 _4673_/D sky130_fd_sc_hd__a22o_1
X_2512_ _4131_/A vssd1 vssd1 vccd1 vccd1 _2512_/X sky130_fd_sc_hd__buf_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3492_ _4703_/Q _3486_/X _4245_/X _3488_/X vssd1 vssd1 vccd1 vccd1 _4703_/D sky130_fd_sc_hd__a22o_1
X_2443_ _2443_/A _2443_/B _2443_/C _2443_/D vssd1 vssd1 vccd1 vccd1 _2443_/Y sky130_fd_sc_hd__nor4_1
X_2374_ input1/X vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__inv_2
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4113_ _4114_/B vssd1 vssd1 vccd1 vccd1 _4113_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2449__B1 _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4044_ _4044_/A vssd1 vssd1 vccd1 vccd1 _4044_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3661__A2 _3633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3949__B1 _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3828_ _3828_/A vssd1 vssd1 vccd1 vccd1 _4505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2924__A1 _4470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3759_ _4556_/Q _3757_/X input8/X _3758_/X vssd1 vssd1 vccd1 vccd1 _4556_/D sky130_fd_sc_hd__a22o_1
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3652__A2 _3647_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2915__A1 _4467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2992_ _4187_/X _2992_/B vssd1 vssd1 vccd1 vccd1 _2992_/X sky130_fd_sc_hd__or2_1
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4731_ _4732_/CLK _4731_/D vssd1 vssd1 vccd1 vccd1 _4731_/Q sky130_fd_sc_hd__dfxtp_1
X_4662_ _4733_/CLK _4662_/D vssd1 vssd1 vccd1 vccd1 _4662_/Q sky130_fd_sc_hd__dfxtp_1
X_3613_ _3328_/A _4650_/Q _3613_/S vssd1 vssd1 vccd1 vccd1 _3614_/A sky130_fd_sc_hd__mux2_1
X_4593_ _4637_/CLK _4593_/D vssd1 vssd1 vccd1 vccd1 _4593_/Q sky130_fd_sc_hd__dfxtp_2
X_3544_ _4213_/X _4679_/Q _3548_/S vssd1 vssd1 vccd1 vccd1 _3545_/A sky130_fd_sc_hd__mux2_1
X_3475_ _3475_/A vssd1 vssd1 vccd1 vccd1 _4711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2426_ _2426_/A _2426_/B vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__or2_1
XFILLER_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2357_ _2355_/A _2355_/B _2355_/Y vssd1 vssd1 vccd1 vccd1 _2357_/Y sky130_fd_sc_hd__a21oi_1
X_2288_ _2288_/A _2288_/B vssd1 vssd1 vccd1 vccd1 _2288_/X sky130_fd_sc_hd__or2_1
X_4027_ input1/X _4037_/B _4029_/C vssd1 vssd1 vccd1 vccd1 _4027_/Y sky130_fd_sc_hd__nor3_1
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2842__B1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4084__B _4092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4304__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3619__A _3655_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4214__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4433__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output88_A _4532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3260_/A _3260_/B vssd1 vssd1 vccd1 vccd1 _3263_/C sky130_fd_sc_hd__nand2_1
XFILLER_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3191_ _3181_/A _3181_/B _3192_/A _3192_/B vssd1 vssd1 vccd1 vccd1 _3193_/C sky130_fd_sc_hd__a22o_1
XFILLER_78_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _2211_/A vssd1 vssd1 vccd1 vccd1 _3962_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4185__A _4769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2975_ _3156_/A _2975_/B vssd1 vssd1 vccd1 vccd1 _2975_/X sky130_fd_sc_hd__or2_1
X_4714_ _4735_/CLK _4714_/D vssd1 vssd1 vccd1 vccd1 _4714_/Q sky130_fd_sc_hd__dfxtp_1
X_4645_ _4649_/CLK _4645_/D vssd1 vssd1 vccd1 vccd1 _4645_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4424__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4576_ _4769_/CLK _4576_/D vssd1 vssd1 vccd1 vccd1 _4576_/Q sky130_fd_sc_hd__dfxtp_1
X_3527_ _3527_/A vssd1 vssd1 vccd1 vccd1 _4687_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3304__A1 _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3458_ _4284_/X _4718_/Q _3458_/S vssd1 vssd1 vccd1 vccd1 _3459_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4079__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2409_ _2409_/A vssd1 vssd1 vccd1 vccd1 _2409_/X sky130_fd_sc_hd__clkbuf_2
X_3389_ _4750_/Q _3374_/A _4254_/X _3375_/A vssd1 vssd1 vccd1 vccd1 _4750_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_48_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3240__B1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2594__A2 _2493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3791__B2 _3786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3791__A1 _4532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4415__S0 _4196_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3349__A _4367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2760_ _2753_/A _2753_/B _2753_/Y vssd1 vssd1 vccd1 vccd1 _2761_/B sky130_fd_sc_hd__a21o_1
XANTENNA__3782__B2 _3303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3782__A1 _4538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2691_ _2702_/B _2691_/B vssd1 vssd1 vccd1 vccd1 _2697_/B sky130_fd_sc_hd__or2_1
XANTENNA__4406__S0 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _4744_/Q _4726_/Q _4693_/Q _4437_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4430_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4139_/X _4134_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4361_/X sky130_fd_sc_hd__mux2_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _4291_/X input39/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4292_/X sky130_fd_sc_hd__mux2_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _4764_/Q _3321_/B vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__nand2_1
XFILLER_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3243_ _2507_/A _3069_/A _2472_/A _3076_/A _3242_/X vssd1 vssd1 vccd1 vccd1 _3244_/D
+ sky130_fd_sc_hd__o221ai_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3174_ _4187_/X _3176_/B vssd1 vssd1 vccd1 vccd1 _3174_/X sky130_fd_sc_hd__and2_1
XFILLER_66_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3222__B1 _3213_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2958_ _2950_/A _2950_/B _2951_/B vssd1 vssd1 vccd1 vccd1 _2959_/A sky130_fd_sc_hd__a21bo_1
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2576__A2 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2889_ _4761_/Q _2889_/B vssd1 vssd1 vccd1 vccd1 _3043_/A sky130_fd_sc_hd__nand2_1
X_4628_ _4629_/CLK _4628_/D vssd1 vssd1 vccd1 vccd1 _4628_/Q sky130_fd_sc_hd__dfxtp_2
X_4559_ _4637_/CLK _4559_/D vssd1 vssd1 vccd1 vccd1 _4559_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_opt_4_0_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_0_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3868__S _3874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2801__A _4470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput72 _4517_/Q vssd1 vssd1 vccd1 vccd1 addr_out[10] sky130_fd_sc_hd__buf_2
Xoutput83 _4527_/Q vssd1 vssd1 vccd1 vccd1 addr_out[20] sky130_fd_sc_hd__buf_2
Xoutput94 _4537_/Q vssd1 vssd1 vccd1 vccd1 addr_out[30] sky130_fd_sc_hd__buf_2
XANTENNA__3819__A2 _3816_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _3944_/A vssd1 vssd1 vccd1 vccd1 _3930_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3861_ _4320_/X _4491_/Q _3863_/S vssd1 vssd1 vccd1 vccd1 _3862_/A sky130_fd_sc_hd__mux2_1
X_3792_ _4531_/Q _3788_/X _4402_/X _3786_/X vssd1 vssd1 vccd1 vccd1 _4531_/D sky130_fd_sc_hd__a22o_1
X_2812_ _2545_/A _2913_/A _2815_/A _2913_/B vssd1 vssd1 vccd1 vccd1 _2819_/A sky130_fd_sc_hd__a22o_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2743_ _2377_/Y _2741_/Y _4194_/X _2742_/B _2742_/Y vssd1 vssd1 vccd1 vccd1 _2743_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3807__A _3814_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2674_ _2674_/A _2679_/A _2679_/B vssd1 vssd1 vccd1 vccd1 _2676_/B sky130_fd_sc_hd__or3_1
XFILLER_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4413_ _4760_/Q _4710_/Q _4677_/Q _4614_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4413_/X sky130_fd_sc_hd__mux4_2
XFILLER_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4344_ _4171_/X _4152_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4344_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4275_ _4029_/Y input48/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4275_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3226_ _2448_/A _4562_/Q _2824_/A _3079_/A vssd1 vssd1 vccd1 vccd1 _3226_/X sky130_fd_sc_hd__o22a_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3691__B1 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3157_ _3152_/A _3152_/B _3152_/Y vssd1 vssd1 vccd1 vccd1 _3157_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3088_ _4567_/Q vssd1 vssd1 vccd1 vccd1 _3089_/A sky130_fd_sc_hd__inv_2
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4092__B _4092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3717__A _3717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4312__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2485__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3627__A _3634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4222__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4162__A1 _2532_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2390_ _2390_/A vssd1 vssd1 vccd1 vccd1 _2390_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4060_ _4060_/A vssd1 vssd1 vccd1 vccd1 _4060_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3011_ _3039_/A _2993_/X _3041_/A _3009_/A _3010_/Y vssd1 vssd1 vccd1 vccd1 _3011_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3913_ _4468_/Q _3906_/X _2543_/A _3909_/X vssd1 vssd1 vccd1 vccd1 _4468_/D sky130_fd_sc_hd__a22o_1
XFILLER_32_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3844_ _4304_/X _4499_/Q _3852_/S vssd1 vssd1 vccd1 vccd1 _3845_/A sky130_fd_sc_hd__mux2_1
X_3775_ _4544_/Q _3771_/X _2500_/A _3772_/X vssd1 vssd1 vccd1 vccd1 _4544_/D sky130_fd_sc_hd__a22o_1
X_2726_ _4631_/Q _2725_/Y _2722_/B vssd1 vssd1 vccd1 vccd1 _2727_/B sky130_fd_sc_hd__o21ai_1
X_2657_ _2721_/A _2721_/B _2657_/C _2725_/B vssd1 vssd1 vccd1 vccd1 _2702_/B sky130_fd_sc_hd__or4_4
X_2588_ _2654_/A _2507_/A _2655_/A _2472_/A _2587_/X vssd1 vssd1 vccd1 vccd1 _2589_/D
+ sky130_fd_sc_hd__o221ai_4
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4327_ _4074_/X _4419_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4327_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4258_ _4257_/X _3981_/A _4354_/S vssd1 vssd1 vccd1 vccd1 _4258_/X sky130_fd_sc_hd__mux2_2
XFILLER_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3209_ _3210_/B _3209_/B _3209_/C _3212_/A vssd1 vssd1 vccd1 vccd1 _3225_/C sky130_fd_sc_hd__or4_2
XFILLER_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4189_ _3968_/Y _3971_/Y _4195_/S vssd1 vssd1 vccd1 vccd1 _4189_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4307__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4144__A1 _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3881__S _3885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2458__B2 _4594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4217__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2630__B2 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3560_ _3560_/A vssd1 vssd1 vccd1 vccd1 _3560_/X sky130_fd_sc_hd__clkbuf_2
X_2511_ input2/X vssd1 vssd1 vccd1 vccd1 _4131_/A sky130_fd_sc_hd__inv_2
X_3491_ _4704_/Q _3486_/X _4241_/X _3488_/X vssd1 vssd1 vccd1 vccd1 _4704_/D sky130_fd_sc_hd__a22o_1
X_2442_ _2373_/A _2377_/A _2379_/X _2441_/X vssd1 vssd1 vccd1 vccd1 _2443_/B sky130_fd_sc_hd__o211ai_2
XFILLER_69_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2373_ _2373_/A vssd1 vssd1 vccd1 vccd1 _2373_/Y sky130_fd_sc_hd__inv_2
X_4112_ _3380_/A input1/X _2493_/A vssd1 vssd1 vccd1 vccd1 _4114_/B sky130_fd_sc_hd__o21ai_1
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4043_ _4375_/X _4250_/S vssd1 vssd1 vccd1 vccd1 _4044_/A sky130_fd_sc_hd__and2_1
XFILLER_17_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3646__B1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3827_ _4280_/X _4505_/Q _3958_/S vssd1 vssd1 vccd1 vccd1 _3828_/A sky130_fd_sc_hd__mux2_1
X_3758_ _3772_/A vssd1 vssd1 vccd1 vccd1 _3758_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2709_ _2709_/A _2709_/B _2709_/C _2708_/X vssd1 vssd1 vccd1 vccd1 _2789_/C sky130_fd_sc_hd__or4b_1
X_3689_ _3696_/A vssd1 vssd1 vccd1 vccd1 _3689_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3637__B1 _2455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3905__A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3628__B1 _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3640__A _3654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2991_ _4192_/X _2991_/B vssd1 vssd1 vccd1 vccd1 _2991_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4730_ _4752_/CLK _4730_/D vssd1 vssd1 vccd1 vccd1 _4730_/Q sky130_fd_sc_hd__dfxtp_1
X_4661_ _4737_/CLK _4661_/D vssd1 vssd1 vccd1 vccd1 _4661_/Q sky130_fd_sc_hd__dfxtp_2
X_3612_ _2211_/A _3320_/A _4205_/X _3330_/Y vssd1 vssd1 vccd1 vccd1 _3613_/S sky130_fd_sc_hd__a211o_1
X_4592_ _4738_/CLK _4592_/D vssd1 vssd1 vccd1 vccd1 _4592_/Q sky130_fd_sc_hd__dfxtp_2
X_3543_ _3543_/A vssd1 vssd1 vccd1 vccd1 _4680_/D sky130_fd_sc_hd__clkbuf_1
X_3474_ _4215_/X _4711_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3475_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2425_ _2426_/A _2426_/B _2417_/X _2419_/X vssd1 vssd1 vccd1 vccd1 _2427_/C sky130_fd_sc_hd__a22o_1
XFILLER_69_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2356_ _4588_/Q _2355_/Y _2254_/B vssd1 vssd1 vccd1 vccd1 _2356_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2287_ _4605_/Q vssd1 vssd1 vccd1 vccd1 _2288_/A sky130_fd_sc_hd__inv_2
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4026_ input1/X _4036_/B _4026_/C vssd1 vssd1 vccd1 vccd1 _4026_/Y sky130_fd_sc_hd__nor3_1
XFILLER_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2842__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4347__A1 _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4320__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4433__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4230__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _3965_/A vssd1 vssd1 vccd1 vccd1 _2211_/A sky130_fd_sc_hd__inv_2
X_3190_ _3179_/A _3179_/B _3179_/Y vssd1 vssd1 vccd1 vccd1 _3192_/B sky130_fd_sc_hd__a21o_1
XFILLER_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2974_ _2968_/A _2968_/B _2968_/Y vssd1 vssd1 vccd1 vccd1 _2975_/B sky130_fd_sc_hd__a21o_1
X_4713_ _4734_/CLK _4713_/D vssd1 vssd1 vccd1 vccd1 _4713_/Q sky130_fd_sc_hd__dfxtp_1
X_4644_ _4644_/CLK _4644_/D vssd1 vssd1 vccd1 vccd1 _4644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4575_ _4769_/CLK _4575_/D vssd1 vssd1 vccd1 vccd1 _4575_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4424__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3526_ _4280_/X _4687_/Q _3530_/S vssd1 vssd1 vccd1 vccd1 _3527_/A sky130_fd_sc_hd__mux2_1
X_3457_ _3457_/A vssd1 vssd1 vccd1 vccd1 _4719_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3304__A2 _4769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2408_ _4365_/X vssd1 vssd1 vccd1 vccd1 _2409_/A sky130_fd_sc_hd__clkinv_2
X_3388_ _4751_/Q _3373_/X _4249_/X _3375_/X vssd1 vssd1 vccd1 vccd1 _4751_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2339_ _4362_/X vssd1 vssd1 vccd1 vccd1 _2340_/A sky130_fd_sc_hd__inv_2
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4095__B _4103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4009_ _4014_/A vssd1 vssd1 vccd1 vccd1 _4013_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4315__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3240__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3791__A2 _3788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4415__S1 _4190_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input32_A addr_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4225__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3782__A2 _3508_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2690_ _2690_/A _2690_/B _2690_/C _2690_/D vssd1 vssd1 vccd1 vccd1 _2789_/A sky130_fd_sc_hd__or4_2
XFILLER_8_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4406__S1 _4202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4360_ _4141_/X _4132_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4360_/X sky130_fd_sc_hd__mux2_1
X_3311_ _2202_/A _3310_/B _4765_/Q _3325_/B vssd1 vssd1 vccd1 vccd1 _3321_/B sky130_fd_sc_hd__o22a_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4020_/Y input39/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4291_/X sky130_fd_sc_hd__mux2_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ input5/X _3242_/B vssd1 vssd1 vccd1 vccd1 _3242_/X sky130_fd_sc_hd__or2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3173_ _3161_/A _3161_/B _3161_/Y vssd1 vssd1 vccd1 vccd1 _3176_/B sky130_fd_sc_hd__a21oi_1
XFILLER_79_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _4755_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2444__A _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2957_ _2951_/A _2951_/B _2951_/Y vssd1 vssd1 vccd1 vccd1 _2957_/Y sky130_fd_sc_hd__a21oi_1
X_2888_ _2805_/X _2809_/X _2819_/Y _2881_/X _2887_/X vssd1 vssd1 vccd1 vccd1 _2889_/B
+ sky130_fd_sc_hd__a41o_2
X_4627_ _4629_/CLK _4627_/D vssd1 vssd1 vccd1 vccd1 _4627_/Q sky130_fd_sc_hd__dfxtp_2
X_4558_ _4558_/CLK _4558_/D vssd1 vssd1 vccd1 vccd1 _4558_/Q sky130_fd_sc_hd__dfxtp_2
X_3509_ _4695_/Q _3508_/X _4411_/X _3303_/X vssd1 vssd1 vccd1 vccd1 _4695_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4489_ _4719_/CLK _4489_/D vssd1 vssd1 vccd1 vccd1 _4489_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4760_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput73 _4518_/Q vssd1 vssd1 vccd1 vccd1 addr_out[11] sky130_fd_sc_hd__buf_2
Xoutput84 _4528_/Q vssd1 vssd1 vccd1 vccd1 addr_out[21] sky130_fd_sc_hd__buf_2
Xoutput95 _4538_/Q vssd1 vssd1 vccd1 vccd1 addr_out[31] sky130_fd_sc_hd__buf_2
XFILLER_95_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_28_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _4747_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _3860_/A vssd1 vssd1 vccd1 vccd1 _4492_/D sky130_fd_sc_hd__clkbuf_1
X_2811_ _4466_/Q vssd1 vssd1 vccd1 vccd1 _2913_/B sky130_fd_sc_hd__inv_2
X_3791_ _4532_/Q _3788_/X _4403_/X _3786_/X vssd1 vssd1 vccd1 vccd1 _4532_/D sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_32_clk_A clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2742_ _4194_/X _2742_/B vssd1 vssd1 vccd1 vccd1 _2742_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2673_ _3092_/A _2670_/B _2277_/Y _2672_/Y vssd1 vssd1 vccd1 vccd1 _2690_/C sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_47_clk_A clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4412_ _4759_/Q _4709_/Q _4676_/Q _4653_/Q _4196_/X _4190_/X vssd1 vssd1 vccd1 vccd1
+ _4412_/X sky130_fd_sc_hd__mux4_1
X_4343_ _4182_/X _4145_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4343_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4274_ _4273_/X input49/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4274_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3225_ _3225_/A _3225_/B _3225_/C _3225_/D vssd1 vssd1 vccd1 vccd1 _3225_/Y sky130_fd_sc_hd__nor4_1
XFILLER_100_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3156_ _3156_/A _3156_/B vssd1 vssd1 vccd1 vccd1 _3156_/X sky130_fd_sc_hd__or2_1
XFILLER_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4571_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3087_ _2266_/X _3086_/X _4352_/X _3084_/Y vssd1 vssd1 vccd1 vccd1 _3087_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _3989_/A vssd1 vssd1 vccd1 vccd1 _4035_/B sky130_fd_sc_hd__clkinv_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3733__A _3771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3879__S _3885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3908__A _3944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3010_ _3008_/X _3002_/A _3004_/X _3009_/C vssd1 vssd1 vccd1 vccd1 _3010_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_49_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3912_ _4469_/Q _3906_/X _2803_/A _3909_/X vssd1 vssd1 vccd1 vccd1 _4469_/D sky130_fd_sc_hd__a22o_1
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3843_ _3900_/S vssd1 vssd1 vccd1 vccd1 _3852_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_20_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_3_0_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_clk/X
+ sky130_fd_sc_hd__clkbuf_16
X_3774_ _4545_/Q _3771_/X _2498_/A _3772_/X vssd1 vssd1 vccd1 vccd1 _4545_/D sky130_fd_sc_hd__a22o_1
X_2725_ _2725_/A _2725_/B vssd1 vssd1 vccd1 vccd1 _2725_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_8_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4626_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2656_ _2656_/A _2770_/A _2768_/A _2768_/B vssd1 vssd1 vccd1 vccd1 _2725_/B sky130_fd_sc_hd__or4_2
X_2587_ _2721_/A input5/X vssd1 vssd1 vccd1 vccd1 _2587_/X sky130_fd_sc_hd__or2_2
X_4326_ _4325_/X _4420_/X _4338_/S vssd1 vssd1 vccd1 vccd1 _4326_/X sky130_fd_sc_hd__mux2_1
X_4257_ _3984_/X _3981_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _4257_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4188_ _4124_/X _2499_/X _4367_/S vssd1 vssd1 vccd1 vccd1 _4188_/X sky130_fd_sc_hd__mux2_1
X_3208_ _3208_/A _3208_/B _3208_/C _3208_/D vssd1 vssd1 vccd1 vccd1 _3212_/A sky130_fd_sc_hd__or4_1
X_3139_ _3136_/Y _3138_/X _2327_/X _3131_/X vssd1 vssd1 vccd1 vccd1 _3143_/B sky130_fd_sc_hd__a22o_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4323__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2458__A2 _4595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output101_A _4515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2630__A2 _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4233__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2510_ _2503_/X _2504_/X _2509_/X vssd1 vssd1 vccd1 vccd1 _2510_/X sky130_fd_sc_hd__a21bo_2
X_3490_ _4705_/Q _3486_/X _4237_/X _3488_/X vssd1 vssd1 vccd1 vccd1 _4705_/D sky130_fd_sc_hd__a22o_1
X_2441_ _2367_/Y _2382_/X _2441_/C _2441_/D vssd1 vssd1 vccd1 vccd1 _2441_/X sky130_fd_sc_hd__and4bb_1
X_2372_ _2244_/Y _2368_/Y _2370_/X vssd1 vssd1 vccd1 vccd1 _2373_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__3894__A1 _4476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4111_ _3381_/D _4013_/A _3380_/A input1/X vssd1 vssd1 vccd1 vccd1 _4111_/X sky130_fd_sc_hd__a22o_1
XFILLER_68_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4042_ _4042_/A vssd1 vssd1 vccd1 vccd1 _4042_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2452__A _2452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3826_ _3826_/A vssd1 vssd1 vccd1 vccd1 _4506_/D sky130_fd_sc_hd__clkbuf_1
X_3757_ _3771_/A vssd1 vssd1 vccd1 vccd1 _3757_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2924__A3 _4471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2708_ _2340_/X _2695_/X _4210_/X _2698_/Y vssd1 vssd1 vccd1 vccd1 _2708_/X sky130_fd_sc_hd__o22a_1
X_3688_ _4602_/Q _3680_/X _2545_/A _3683_/X vssd1 vssd1 vccd1 vccd1 _4602_/D sky130_fd_sc_hd__a22o_1
X_2639_ _2636_/A _2638_/X _2636_/C vssd1 vssd1 vccd1 vccd1 _2639_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__3885__A1 _4480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4309_ _4093_/X _4427_/X _4337_/S vssd1 vssd1 vccd1 vccd1 _4309_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3637__A1 _4637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4318__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3892__S _3896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2376__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input62_A data_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2537__A _2537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4228__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2990_ _4187_/X _2992_/B vssd1 vssd1 vccd1 vccd1 _3039_/B sky130_fd_sc_hd__and2_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4733_/CLK _4660_/D vssd1 vssd1 vccd1 vccd1 _4660_/Q sky130_fd_sc_hd__dfxtp_1
X_3611_ _3611_/A vssd1 vssd1 vccd1 vccd1 _4651_/D sky130_fd_sc_hd__clkbuf_1
X_4591_ _4634_/CLK _4591_/D vssd1 vssd1 vccd1 vccd1 _4591_/Q sky130_fd_sc_hd__dfxtp_2
X_3542_ _4340_/X _4680_/Q _3548_/S vssd1 vssd1 vccd1 vccd1 _3543_/A sky130_fd_sc_hd__mux2_1
X_3473_ _3473_/A vssd1 vssd1 vccd1 vccd1 _4712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2424_ _2471_/B _2418_/X _2355_/B vssd1 vssd1 vccd1 vccd1 _2426_/B sky130_fd_sc_hd__a21bo_1
X_2355_ _2355_/A _2355_/B vssd1 vssd1 vccd1 vccd1 _2355_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2286_ _4606_/Q vssd1 vssd1 vccd1 vccd1 _2286_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2447__A _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4025_ input1/X _4035_/B _4026_/C vssd1 vssd1 vccd1 vccd1 _4025_/Y sky130_fd_sc_hd__nor3_1
XFILLER_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3809_ _3816_/A vssd1 vssd1 vccd1 vccd1 _3809_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4283__A1 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3916__A _3923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__4274__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2973_ _3154_/A _2973_/B vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__or2_1
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2588__B2 _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4712_ _4733_/CLK _4712_/D vssd1 vssd1 vccd1 vccd1 _4712_/Q sky130_fd_sc_hd__dfxtp_1
X_4643_ _4644_/CLK _4643_/D vssd1 vssd1 vccd1 vccd1 _4643_/Q sky130_fd_sc_hd__dfxtp_1
X_4574_ _4738_/CLK _4574_/D vssd1 vssd1 vccd1 vccd1 _4574_/Q sky130_fd_sc_hd__dfxtp_1
X_3525_ _3525_/A vssd1 vssd1 vccd1 vccd1 _4688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3456_ _4282_/X _4719_/Q _3458_/S vssd1 vssd1 vccd1 vccd1 _3457_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2407_ _2407_/A _2407_/B _2407_/C _2407_/D vssd1 vssd1 vccd1 vccd1 _2430_/A sky130_fd_sc_hd__or4_1
X_3387_ _3387_/A vssd1 vssd1 vccd1 vccd1 _4752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2338_ _4210_/X _2337_/X _2327_/X _2329_/Y vssd1 vssd1 vccd1 vccd1 _2344_/B sky130_fd_sc_hd__a22o_1
X_2269_ _4191_/X vssd1 vssd1 vccd1 vccd1 _2916_/A sky130_fd_sc_hd__inv_2
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4008_ _4008_/A vssd1 vssd1 vccd1 vccd1 _4008_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4265__A1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3776__B1 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2579__B2 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3736__A _3772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4331__S _4337_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3700__B1 _2455_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_A addr_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4256__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2815__A _2815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3767__B1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4241__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output93_A _4509_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3310_ _4338_/S _3310_/B vssd1 vssd1 vccd1 vccd1 _3319_/A sky130_fd_sc_hd__or2_1
XFILLER_98_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ _4289_/X input40/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4290_/X sky130_fd_sc_hd__mux2_1
X_3241_ _4136_/A _4555_/Q _2484_/A _4554_/Q _3240_/X vssd1 vssd1 vccd1 vccd1 _3244_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3381__A _3965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3172_ _4194_/X _3170_/B _3171_/X vssd1 vssd1 vccd1 vccd1 _3172_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_6_clk_A clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4247__A1 _4375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2956_ _2956_/A _2956_/B _2956_/C _2955_/X vssd1 vssd1 vccd1 vccd1 _3032_/C sky130_fd_sc_hd__or4b_1
XFILLER_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2887_ _2535_/A _2806_/Y _2882_/Y _2886_/X vssd1 vssd1 vccd1 vccd1 _2887_/X sky130_fd_sc_hd__o22a_1
X_4626_ _4626_/CLK _4626_/D vssd1 vssd1 vccd1 vccd1 _4626_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3556__A _4354_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4557_ _4558_/CLK _4557_/D vssd1 vssd1 vccd1 vccd1 _4557_/Q sky130_fd_sc_hd__dfxtp_2
X_3508_ _3788_/A vssd1 vssd1 vccd1 vccd1 _3508_/X sky130_fd_sc_hd__buf_2
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4488_ _4760_/CLK _4488_/D vssd1 vssd1 vccd1 vccd1 _4488_/Q sky130_fd_sc_hd__dfxtp_4
X_3439_ _3439_/A vssd1 vssd1 vccd1 vccd1 _4727_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2497__B1 _2492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4326__S _4338_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3749__B1 _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2370__A _4665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3466__A _3484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3921__B1 _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput85 _4529_/Q vssd1 vssd1 vccd1 vccd1 addr_out[22] sky130_fd_sc_hd__buf_2
XFILLER_95_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput74 _4519_/Q vssd1 vssd1 vccd1 vccd1 addr_out[12] sky130_fd_sc_hd__buf_2
XANTENNA__2488__B1 _2472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput96 _4510_/Q vssd1 vssd1 vccd1 vccd1 addr_out[3] sky130_fd_sc_hd__buf_2
XFILLER_88_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output131_A _4479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4229__A1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2545__A _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4236__S _4339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2810_ _4467_/Q vssd1 vssd1 vccd1 vccd1 _2913_/A sky130_fd_sc_hd__inv_2
X_3790_ _4533_/Q _3788_/X _4404_/X _3786_/X vssd1 vssd1 vccd1 vccd1 _4533_/D sky130_fd_sc_hd__a22o_1
XANTENNA__4401__A1 _4598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2741_ _2741_/A vssd1 vssd1 vccd1 vccd1 _2741_/Y sky130_fd_sc_hd__inv_2
X_4411_ _4700_/Q _4665_/Q _4663_/Q _4661_/Q _4203_/X _4202_/X vssd1 vssd1 vccd1 vccd1
+ _4411_/X sky130_fd_sc_hd__mux4_1
X_2672_ _2672_/A vssd1 vssd1 vccd1 vccd1 _2672_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3912__B1 _2803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4342_ _4169_/Y _2816_/A _4367_/S vssd1 vssd1 vccd1 vccd1 _4342_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4273_ _4032_/Y input49/X _4339_/S vssd1 vssd1 vccd1 vccd1 _4273_/X sky130_fd_sc_hd__mux2_1
X_3224_ _2377_/A _3169_/A _3171_/X _3223_/X vssd1 vssd1 vccd1 vccd1 _3225_/B sky130_fd_sc_hd__o211ai_1
.ends

