VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 1496.000 7.270 1500.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.690 1496.000 1315.970 1500.000 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1243.080 1500.000 1243.680 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1287.960 4.000 1288.560 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.330 0.000 1239.610 4.000 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.030 0.000 1260.310 4.000 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1283.880 1500.000 1284.480 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.890 0.000 1302.170 4.000 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.920 4.000 1303.520 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.130 1496.000 1345.410 1500.000 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.570 1496.000 1374.850 1500.000 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 1496.000 330.650 1500.000 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1345.760 1500.000 1346.360 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1331.480 4.000 1332.080 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1386.560 1500.000 1387.160 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1406.960 1500.000 1407.560 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 1496.000 1404.290 1500.000 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1428.040 1500.000 1428.640 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.720 4.000 1361.320 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 0.000 1406.130 4.000 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 0.000 1426.830 4.000 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.710 0.000 1447.990 4.000 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1419.200 4.000 1419.800 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1433.480 4.000 1434.080 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1448.440 4.000 1449.040 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.170 1496.000 1448.450 1500.000 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.890 1496.000 1463.170 1500.000 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.720 4.000 1463.320 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.330 1496.000 1492.610 1500.000 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1477.680 4.000 1478.280 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 338.680 1500.000 339.280 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 1496.000 389.530 1500.000 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 1496.000 492.570 1500.000 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 400.560 1500.000 401.160 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 1496.000 536.270 1500.000 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.160 4.000 414.760 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1496.000 109.850 1500.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 523.640 1500.000 524.240 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 1496.000 595.150 1500.000 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 1496.000 639.310 1500.000 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.680 4.000 662.280 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 729.000 1500.000 729.600 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 1496.000 727.630 1500.000 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 1496.000 742.350 1500.000 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 1496.000 757.070 1500.000 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 1496.000 771.790 1500.000 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 1496.000 786.510 1500.000 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 811.280 1500.000 811.880 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 831.680 1500.000 832.280 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 1496.000 815.950 1500.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.680 4.000 764.280 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 873.160 1500.000 873.760 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 1496.000 860.110 1500.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 1496.000 183.450 1500.000 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 1496.000 874.830 1500.000 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 1496.000 889.550 1500.000 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.160 4.000 822.760 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 1496.000 904.270 1500.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 934.360 1500.000 934.960 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 4.000 852.000 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.680 4.000 866.280 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 955.440 1500.000 956.040 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 975.840 1500.000 976.440 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 1496.000 963.150 1500.000 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.590 1496.000 977.870 1500.000 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 0.000 885.410 4.000 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.830 0.000 906.110 4.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 996.240 1500.000 996.840 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 953.400 4.000 954.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.530 0.000 926.810 4.000 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 967.680 4.000 968.280 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 1496.000 271.770 1500.000 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.030 1496.000 1007.310 1500.000 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.200 4.000 1011.800 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1055.400 4.000 1056.000 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1078.520 1500.000 1079.120 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1098.920 1500.000 1099.520 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 0.000 1010.530 4.000 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1069.680 4.000 1070.280 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1083.960 4.000 1084.560 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.920 4.000 1099.520 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1113.200 4.000 1113.800 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1140.400 1500.000 1141.000 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.160 4.000 1128.760 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 1496.000 1109.890 1500.000 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.050 1496.000 1139.330 1500.000 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.510 0.000 1093.790 4.000 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.720 4.000 1157.320 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 0.000 1135.190 4.000 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.490 1496.000 1168.770 1500.000 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 1496.000 1183.490 1500.000 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1171.680 4.000 1172.280 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.650 1496.000 1212.930 1500.000 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1215.200 4.000 1215.800 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1201.600 1500.000 1202.200 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 1496.000 1227.650 1500.000 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.470 0.000 1197.750 4.000 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.720 4.000 1259.320 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.530 1496.000 1271.810 1500.000 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.250 1496.000 1286.530 1500.000 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 30.640 1500.000 31.240 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 1496.000 345.370 1500.000 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 1496.000 374.810 1500.000 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 1496.000 404.250 1500.000 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 1496.000 433.690 1500.000 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 379.480 1500.000 380.080 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 420.960 1500.000 421.560 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 1496.000 124.570 1500.000 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 482.840 1500.000 483.440 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 544.040 1500.000 544.640 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 585.520 1500.000 586.120 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1496.000 654.030 1500.000 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.160 4.000 618.760 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 667.800 1500.000 668.400 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 153.720 1500.000 154.320 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1496.000 212.890 1500.000 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 1496.000 286.490 1500.000 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1496.000 315.930 1500.000 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 1496.000 65.690 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 1496.000 95.130 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 10.240 1500.000 10.840 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 1496.000 80.410 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 359.080 1500.000 359.680 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 1496.000 448.410 1500.000 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 133.320 1500.000 133.920 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 174.120 1500.000 174.720 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 1496.000 227.610 1500.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 215.600 1500.000 216.200 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 276.800 1500.000 277.400 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 51.040 1500.000 51.640 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1273.680 4.000 1274.280 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 1496.000 1330.690 1500.000 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 4.000 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1263.480 1500.000 1264.080 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.730 0.000 1281.010 4.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1304.280 1500.000 1304.880 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.590 0.000 1322.870 4.000 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1317.200 4.000 1317.800 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.850 1496.000 1360.130 1500.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1325.360 1500.000 1325.960 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 318.280 1500.000 318.880 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1366.160 1500.000 1366.760 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.290 1496.000 1389.570 1500.000 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1346.440 4.000 1347.040 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.290 0.000 1343.570 4.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 0.000 1364.270 4.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1375.680 4.000 1376.280 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1389.960 4.000 1390.560 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.920 4.000 1405.520 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 1496.000 1419.010 1500.000 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1448.440 1500.000 1449.040 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.450 1496.000 1433.730 1500.000 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1468.840 1500.000 1469.440 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.610 1496.000 1477.890 1500.000 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 0.000 1489.390 4.000 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1489.240 1500.000 1489.840 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.960 4.000 1492.560 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 1496.000 463.130 1500.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 441.360 1500.000 441.960 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 461.760 1500.000 462.360 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 91.840 1500.000 92.440 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 503.240 1500.000 503.840 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 564.440 1500.000 565.040 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 1496.000 580.430 1500.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 1496.000 609.870 1500.000 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 0.000 531.210 4.000 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 605.920 1500.000 606.520 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 1496.000 139.290 1500.000 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 688.200 1500.000 688.800 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 708.600 1500.000 709.200 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 1496.000 712.910 1500.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 749.400 1500.000 750.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 770.480 1500.000 771.080 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 790.880 1500.000 791.480 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 1496.000 154.010 1500.000 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 1496.000 801.230 1500.000 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 1496.000 830.670 1500.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 852.080 1500.000 852.680 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 1496.000 845.390 1500.000 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 893.560 1500.000 894.160 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 1496.000 198.170 1500.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.200 4.000 807.800 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 913.960 1500.000 914.560 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 0.000 780.990 4.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.710 1496.000 918.990 1500.000 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 1496.000 933.710 1500.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 1496.000 948.430 1500.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 1496.000 242.330 1500.000 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.920 4.000 895.520 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 0.000 864.250 4.000 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 1496.000 992.590 1500.000 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.200 4.000 909.800 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.160 4.000 924.760 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1016.640 1500.000 1017.240 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.690 0.000 947.970 4.000 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.960 4.000 982.560 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1037.040 1500.000 1037.640 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 194.520 1500.000 195.120 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 0.000 968.670 4.000 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.160 4.000 1026.760 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 1496.000 1021.570 1500.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1058.120 1500.000 1058.720 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 1496.000 1036.290 1500.000 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.090 0.000 989.370 4.000 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.730 1496.000 1051.010 1500.000 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1119.320 1500.000 1119.920 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 0.000 1031.230 4.000 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 1496.000 1065.730 1500.000 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 1496.000 301.210 1500.000 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.170 1496.000 1080.450 1500.000 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 1496.000 1095.170 1500.000 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 0.000 1051.930 4.000 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1160.800 1500.000 1161.400 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 1496.000 1124.610 1500.000 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.770 1496.000 1154.050 1500.000 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.070 0.000 1156.350 4.000 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1181.200 1500.000 1181.800 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 256.400 1500.000 257.000 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 1496.000 1198.210 1500.000 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1185.960 4.000 1186.560 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.920 4.000 1201.520 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 4.000 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.160 4.000 1230.760 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1244.440 4.000 1245.040 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.090 1496.000 1242.370 1500.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.810 1496.000 1257.090 1500.000 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1222.000 1500.000 1222.600 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.970 1496.000 1301.250 1500.000 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 297.880 1500.000 298.480 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 1496.000 36.250 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 1496.000 50.970 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 71.440 1500.000 72.040 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 1496.000 360.090 1500.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 1496.000 418.970 1500.000 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 1496.000 477.850 1500.000 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 1496.000 507.290 1500.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 1496.000 521.550 1500.000 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1496.000 550.990 1500.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 112.920 1500.000 113.520 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 1496.000 565.710 1500.000 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.160 4.000 516.760 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 0.000 510.510 4.000 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 1496.000 624.590 1500.000 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 626.320 1500.000 626.920 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 1496.000 668.750 1500.000 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 1496.000 683.470 1500.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 646.720 1500.000 647.320 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 1496.000 698.190 1500.000 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 1496.000 168.730 1500.000 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 1496.000 257.050 1500.000 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 236.000 1500.000 236.600 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 1496.000 21.530 1500.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 7.860 1494.080 1488.080 ;
      LAYER met2 ;
        RECT 7.550 1495.720 20.970 1496.410 ;
        RECT 21.810 1495.720 35.690 1496.410 ;
        RECT 36.530 1495.720 50.410 1496.410 ;
        RECT 51.250 1495.720 65.130 1496.410 ;
        RECT 65.970 1495.720 79.850 1496.410 ;
        RECT 80.690 1495.720 94.570 1496.410 ;
        RECT 95.410 1495.720 109.290 1496.410 ;
        RECT 110.130 1495.720 124.010 1496.410 ;
        RECT 124.850 1495.720 138.730 1496.410 ;
        RECT 139.570 1495.720 153.450 1496.410 ;
        RECT 154.290 1495.720 168.170 1496.410 ;
        RECT 169.010 1495.720 182.890 1496.410 ;
        RECT 183.730 1495.720 197.610 1496.410 ;
        RECT 198.450 1495.720 212.330 1496.410 ;
        RECT 213.170 1495.720 227.050 1496.410 ;
        RECT 227.890 1495.720 241.770 1496.410 ;
        RECT 242.610 1495.720 256.490 1496.410 ;
        RECT 257.330 1495.720 271.210 1496.410 ;
        RECT 272.050 1495.720 285.930 1496.410 ;
        RECT 286.770 1495.720 300.650 1496.410 ;
        RECT 301.490 1495.720 315.370 1496.410 ;
        RECT 316.210 1495.720 330.090 1496.410 ;
        RECT 330.930 1495.720 344.810 1496.410 ;
        RECT 345.650 1495.720 359.530 1496.410 ;
        RECT 360.370 1495.720 374.250 1496.410 ;
        RECT 375.090 1495.720 388.970 1496.410 ;
        RECT 389.810 1495.720 403.690 1496.410 ;
        RECT 404.530 1495.720 418.410 1496.410 ;
        RECT 419.250 1495.720 433.130 1496.410 ;
        RECT 433.970 1495.720 447.850 1496.410 ;
        RECT 448.690 1495.720 462.570 1496.410 ;
        RECT 463.410 1495.720 477.290 1496.410 ;
        RECT 478.130 1495.720 492.010 1496.410 ;
        RECT 492.850 1495.720 506.730 1496.410 ;
        RECT 507.570 1495.720 520.990 1496.410 ;
        RECT 521.830 1495.720 535.710 1496.410 ;
        RECT 536.550 1495.720 550.430 1496.410 ;
        RECT 551.270 1495.720 565.150 1496.410 ;
        RECT 565.990 1495.720 579.870 1496.410 ;
        RECT 580.710 1495.720 594.590 1496.410 ;
        RECT 595.430 1495.720 609.310 1496.410 ;
        RECT 610.150 1495.720 624.030 1496.410 ;
        RECT 624.870 1495.720 638.750 1496.410 ;
        RECT 639.590 1495.720 653.470 1496.410 ;
        RECT 654.310 1495.720 668.190 1496.410 ;
        RECT 669.030 1495.720 682.910 1496.410 ;
        RECT 683.750 1495.720 697.630 1496.410 ;
        RECT 698.470 1495.720 712.350 1496.410 ;
        RECT 713.190 1495.720 727.070 1496.410 ;
        RECT 727.910 1495.720 741.790 1496.410 ;
        RECT 742.630 1495.720 756.510 1496.410 ;
        RECT 757.350 1495.720 771.230 1496.410 ;
        RECT 772.070 1495.720 785.950 1496.410 ;
        RECT 786.790 1495.720 800.670 1496.410 ;
        RECT 801.510 1495.720 815.390 1496.410 ;
        RECT 816.230 1495.720 830.110 1496.410 ;
        RECT 830.950 1495.720 844.830 1496.410 ;
        RECT 845.670 1495.720 859.550 1496.410 ;
        RECT 860.390 1495.720 874.270 1496.410 ;
        RECT 875.110 1495.720 888.990 1496.410 ;
        RECT 889.830 1495.720 903.710 1496.410 ;
        RECT 904.550 1495.720 918.430 1496.410 ;
        RECT 919.270 1495.720 933.150 1496.410 ;
        RECT 933.990 1495.720 947.870 1496.410 ;
        RECT 948.710 1495.720 962.590 1496.410 ;
        RECT 963.430 1495.720 977.310 1496.410 ;
        RECT 978.150 1495.720 992.030 1496.410 ;
        RECT 992.870 1495.720 1006.750 1496.410 ;
        RECT 1007.590 1495.720 1021.010 1496.410 ;
        RECT 1021.850 1495.720 1035.730 1496.410 ;
        RECT 1036.570 1495.720 1050.450 1496.410 ;
        RECT 1051.290 1495.720 1065.170 1496.410 ;
        RECT 1066.010 1495.720 1079.890 1496.410 ;
        RECT 1080.730 1495.720 1094.610 1496.410 ;
        RECT 1095.450 1495.720 1109.330 1496.410 ;
        RECT 1110.170 1495.720 1124.050 1496.410 ;
        RECT 1124.890 1495.720 1138.770 1496.410 ;
        RECT 1139.610 1495.720 1153.490 1496.410 ;
        RECT 1154.330 1495.720 1168.210 1496.410 ;
        RECT 1169.050 1495.720 1182.930 1496.410 ;
        RECT 1183.770 1495.720 1197.650 1496.410 ;
        RECT 1198.490 1495.720 1212.370 1496.410 ;
        RECT 1213.210 1495.720 1227.090 1496.410 ;
        RECT 1227.930 1495.720 1241.810 1496.410 ;
        RECT 1242.650 1495.720 1256.530 1496.410 ;
        RECT 1257.370 1495.720 1271.250 1496.410 ;
        RECT 1272.090 1495.720 1285.970 1496.410 ;
        RECT 1286.810 1495.720 1300.690 1496.410 ;
        RECT 1301.530 1495.720 1315.410 1496.410 ;
        RECT 1316.250 1495.720 1330.130 1496.410 ;
        RECT 1330.970 1495.720 1344.850 1496.410 ;
        RECT 1345.690 1495.720 1359.570 1496.410 ;
        RECT 1360.410 1495.720 1374.290 1496.410 ;
        RECT 1375.130 1495.720 1389.010 1496.410 ;
        RECT 1389.850 1495.720 1403.730 1496.410 ;
        RECT 1404.570 1495.720 1418.450 1496.410 ;
        RECT 1419.290 1495.720 1433.170 1496.410 ;
        RECT 1434.010 1495.720 1447.890 1496.410 ;
        RECT 1448.730 1495.720 1462.610 1496.410 ;
        RECT 1463.450 1495.720 1477.330 1496.410 ;
        RECT 1478.170 1495.720 1492.050 1496.410 ;
        RECT 6.990 4.280 1492.540 1495.720 ;
        RECT 6.990 3.670 9.930 4.280 ;
        RECT 10.770 3.670 30.630 4.280 ;
        RECT 31.470 3.670 51.330 4.280 ;
        RECT 52.170 3.670 72.030 4.280 ;
        RECT 72.870 3.670 93.190 4.280 ;
        RECT 94.030 3.670 113.890 4.280 ;
        RECT 114.730 3.670 134.590 4.280 ;
        RECT 135.430 3.670 155.750 4.280 ;
        RECT 156.590 3.670 176.450 4.280 ;
        RECT 177.290 3.670 197.150 4.280 ;
        RECT 197.990 3.670 217.850 4.280 ;
        RECT 218.690 3.670 239.010 4.280 ;
        RECT 239.850 3.670 259.710 4.280 ;
        RECT 260.550 3.670 280.410 4.280 ;
        RECT 281.250 3.670 301.570 4.280 ;
        RECT 302.410 3.670 322.270 4.280 ;
        RECT 323.110 3.670 342.970 4.280 ;
        RECT 343.810 3.670 363.670 4.280 ;
        RECT 364.510 3.670 384.830 4.280 ;
        RECT 385.670 3.670 405.530 4.280 ;
        RECT 406.370 3.670 426.230 4.280 ;
        RECT 427.070 3.670 447.390 4.280 ;
        RECT 448.230 3.670 468.090 4.280 ;
        RECT 468.930 3.670 488.790 4.280 ;
        RECT 489.630 3.670 509.950 4.280 ;
        RECT 510.790 3.670 530.650 4.280 ;
        RECT 531.490 3.670 551.350 4.280 ;
        RECT 552.190 3.670 572.050 4.280 ;
        RECT 572.890 3.670 593.210 4.280 ;
        RECT 594.050 3.670 613.910 4.280 ;
        RECT 614.750 3.670 634.610 4.280 ;
        RECT 635.450 3.670 655.770 4.280 ;
        RECT 656.610 3.670 676.470 4.280 ;
        RECT 677.310 3.670 697.170 4.280 ;
        RECT 698.010 3.670 717.870 4.280 ;
        RECT 718.710 3.670 739.030 4.280 ;
        RECT 739.870 3.670 759.730 4.280 ;
        RECT 760.570 3.670 780.430 4.280 ;
        RECT 781.270 3.670 801.590 4.280 ;
        RECT 802.430 3.670 822.290 4.280 ;
        RECT 823.130 3.670 842.990 4.280 ;
        RECT 843.830 3.670 863.690 4.280 ;
        RECT 864.530 3.670 884.850 4.280 ;
        RECT 885.690 3.670 905.550 4.280 ;
        RECT 906.390 3.670 926.250 4.280 ;
        RECT 927.090 3.670 947.410 4.280 ;
        RECT 948.250 3.670 968.110 4.280 ;
        RECT 968.950 3.670 988.810 4.280 ;
        RECT 989.650 3.670 1009.970 4.280 ;
        RECT 1010.810 3.670 1030.670 4.280 ;
        RECT 1031.510 3.670 1051.370 4.280 ;
        RECT 1052.210 3.670 1072.070 4.280 ;
        RECT 1072.910 3.670 1093.230 4.280 ;
        RECT 1094.070 3.670 1113.930 4.280 ;
        RECT 1114.770 3.670 1134.630 4.280 ;
        RECT 1135.470 3.670 1155.790 4.280 ;
        RECT 1156.630 3.670 1176.490 4.280 ;
        RECT 1177.330 3.670 1197.190 4.280 ;
        RECT 1198.030 3.670 1217.890 4.280 ;
        RECT 1218.730 3.670 1239.050 4.280 ;
        RECT 1239.890 3.670 1259.750 4.280 ;
        RECT 1260.590 3.670 1280.450 4.280 ;
        RECT 1281.290 3.670 1301.610 4.280 ;
        RECT 1302.450 3.670 1322.310 4.280 ;
        RECT 1323.150 3.670 1343.010 4.280 ;
        RECT 1343.850 3.670 1363.710 4.280 ;
        RECT 1364.550 3.670 1384.870 4.280 ;
        RECT 1385.710 3.670 1405.570 4.280 ;
        RECT 1406.410 3.670 1426.270 4.280 ;
        RECT 1427.110 3.670 1447.430 4.280 ;
        RECT 1448.270 3.670 1468.130 4.280 ;
        RECT 1468.970 3.670 1488.830 4.280 ;
        RECT 1489.670 3.670 1492.540 4.280 ;
      LAYER met3 ;
        RECT 4.400 1491.560 1496.000 1492.425 ;
        RECT 4.000 1490.240 1496.000 1491.560 ;
        RECT 4.000 1488.840 1495.600 1490.240 ;
        RECT 4.000 1478.680 1496.000 1488.840 ;
        RECT 4.400 1477.280 1496.000 1478.680 ;
        RECT 4.000 1469.840 1496.000 1477.280 ;
        RECT 4.000 1468.440 1495.600 1469.840 ;
        RECT 4.000 1463.720 1496.000 1468.440 ;
        RECT 4.400 1462.320 1496.000 1463.720 ;
        RECT 4.000 1449.440 1496.000 1462.320 ;
        RECT 4.400 1448.040 1495.600 1449.440 ;
        RECT 4.000 1434.480 1496.000 1448.040 ;
        RECT 4.400 1433.080 1496.000 1434.480 ;
        RECT 4.000 1429.040 1496.000 1433.080 ;
        RECT 4.000 1427.640 1495.600 1429.040 ;
        RECT 4.000 1420.200 1496.000 1427.640 ;
        RECT 4.400 1418.800 1496.000 1420.200 ;
        RECT 4.000 1407.960 1496.000 1418.800 ;
        RECT 4.000 1406.560 1495.600 1407.960 ;
        RECT 4.000 1405.920 1496.000 1406.560 ;
        RECT 4.400 1404.520 1496.000 1405.920 ;
        RECT 4.000 1390.960 1496.000 1404.520 ;
        RECT 4.400 1389.560 1496.000 1390.960 ;
        RECT 4.000 1387.560 1496.000 1389.560 ;
        RECT 4.000 1386.160 1495.600 1387.560 ;
        RECT 4.000 1376.680 1496.000 1386.160 ;
        RECT 4.400 1375.280 1496.000 1376.680 ;
        RECT 4.000 1367.160 1496.000 1375.280 ;
        RECT 4.000 1365.760 1495.600 1367.160 ;
        RECT 4.000 1361.720 1496.000 1365.760 ;
        RECT 4.400 1360.320 1496.000 1361.720 ;
        RECT 4.000 1347.440 1496.000 1360.320 ;
        RECT 4.400 1346.760 1496.000 1347.440 ;
        RECT 4.400 1346.040 1495.600 1346.760 ;
        RECT 4.000 1345.360 1495.600 1346.040 ;
        RECT 4.000 1332.480 1496.000 1345.360 ;
        RECT 4.400 1331.080 1496.000 1332.480 ;
        RECT 4.000 1326.360 1496.000 1331.080 ;
        RECT 4.000 1324.960 1495.600 1326.360 ;
        RECT 4.000 1318.200 1496.000 1324.960 ;
        RECT 4.400 1316.800 1496.000 1318.200 ;
        RECT 4.000 1305.280 1496.000 1316.800 ;
        RECT 4.000 1303.920 1495.600 1305.280 ;
        RECT 4.400 1303.880 1495.600 1303.920 ;
        RECT 4.400 1302.520 1496.000 1303.880 ;
        RECT 4.000 1288.960 1496.000 1302.520 ;
        RECT 4.400 1287.560 1496.000 1288.960 ;
        RECT 4.000 1284.880 1496.000 1287.560 ;
        RECT 4.000 1283.480 1495.600 1284.880 ;
        RECT 4.000 1274.680 1496.000 1283.480 ;
        RECT 4.400 1273.280 1496.000 1274.680 ;
        RECT 4.000 1264.480 1496.000 1273.280 ;
        RECT 4.000 1263.080 1495.600 1264.480 ;
        RECT 4.000 1259.720 1496.000 1263.080 ;
        RECT 4.400 1258.320 1496.000 1259.720 ;
        RECT 4.000 1245.440 1496.000 1258.320 ;
        RECT 4.400 1244.080 1496.000 1245.440 ;
        RECT 4.400 1244.040 1495.600 1244.080 ;
        RECT 4.000 1242.680 1495.600 1244.040 ;
        RECT 4.000 1231.160 1496.000 1242.680 ;
        RECT 4.400 1229.760 1496.000 1231.160 ;
        RECT 4.000 1223.000 1496.000 1229.760 ;
        RECT 4.000 1221.600 1495.600 1223.000 ;
        RECT 4.000 1216.200 1496.000 1221.600 ;
        RECT 4.400 1214.800 1496.000 1216.200 ;
        RECT 4.000 1202.600 1496.000 1214.800 ;
        RECT 4.000 1201.920 1495.600 1202.600 ;
        RECT 4.400 1201.200 1495.600 1201.920 ;
        RECT 4.400 1200.520 1496.000 1201.200 ;
        RECT 4.000 1186.960 1496.000 1200.520 ;
        RECT 4.400 1185.560 1496.000 1186.960 ;
        RECT 4.000 1182.200 1496.000 1185.560 ;
        RECT 4.000 1180.800 1495.600 1182.200 ;
        RECT 4.000 1172.680 1496.000 1180.800 ;
        RECT 4.400 1171.280 1496.000 1172.680 ;
        RECT 4.000 1161.800 1496.000 1171.280 ;
        RECT 4.000 1160.400 1495.600 1161.800 ;
        RECT 4.000 1157.720 1496.000 1160.400 ;
        RECT 4.400 1156.320 1496.000 1157.720 ;
        RECT 4.000 1143.440 1496.000 1156.320 ;
        RECT 4.400 1142.040 1496.000 1143.440 ;
        RECT 4.000 1141.400 1496.000 1142.040 ;
        RECT 4.000 1140.000 1495.600 1141.400 ;
        RECT 4.000 1129.160 1496.000 1140.000 ;
        RECT 4.400 1127.760 1496.000 1129.160 ;
        RECT 4.000 1120.320 1496.000 1127.760 ;
        RECT 4.000 1118.920 1495.600 1120.320 ;
        RECT 4.000 1114.200 1496.000 1118.920 ;
        RECT 4.400 1112.800 1496.000 1114.200 ;
        RECT 4.000 1099.920 1496.000 1112.800 ;
        RECT 4.400 1098.520 1495.600 1099.920 ;
        RECT 4.000 1084.960 1496.000 1098.520 ;
        RECT 4.400 1083.560 1496.000 1084.960 ;
        RECT 4.000 1079.520 1496.000 1083.560 ;
        RECT 4.000 1078.120 1495.600 1079.520 ;
        RECT 4.000 1070.680 1496.000 1078.120 ;
        RECT 4.400 1069.280 1496.000 1070.680 ;
        RECT 4.000 1059.120 1496.000 1069.280 ;
        RECT 4.000 1057.720 1495.600 1059.120 ;
        RECT 4.000 1056.400 1496.000 1057.720 ;
        RECT 4.400 1055.000 1496.000 1056.400 ;
        RECT 4.000 1041.440 1496.000 1055.000 ;
        RECT 4.400 1040.040 1496.000 1041.440 ;
        RECT 4.000 1038.040 1496.000 1040.040 ;
        RECT 4.000 1036.640 1495.600 1038.040 ;
        RECT 4.000 1027.160 1496.000 1036.640 ;
        RECT 4.400 1025.760 1496.000 1027.160 ;
        RECT 4.000 1017.640 1496.000 1025.760 ;
        RECT 4.000 1016.240 1495.600 1017.640 ;
        RECT 4.000 1012.200 1496.000 1016.240 ;
        RECT 4.400 1010.800 1496.000 1012.200 ;
        RECT 4.000 997.920 1496.000 1010.800 ;
        RECT 4.400 997.240 1496.000 997.920 ;
        RECT 4.400 996.520 1495.600 997.240 ;
        RECT 4.000 995.840 1495.600 996.520 ;
        RECT 4.000 982.960 1496.000 995.840 ;
        RECT 4.400 981.560 1496.000 982.960 ;
        RECT 4.000 976.840 1496.000 981.560 ;
        RECT 4.000 975.440 1495.600 976.840 ;
        RECT 4.000 968.680 1496.000 975.440 ;
        RECT 4.400 967.280 1496.000 968.680 ;
        RECT 4.000 956.440 1496.000 967.280 ;
        RECT 4.000 955.040 1495.600 956.440 ;
        RECT 4.000 954.400 1496.000 955.040 ;
        RECT 4.400 953.000 1496.000 954.400 ;
        RECT 4.000 939.440 1496.000 953.000 ;
        RECT 4.400 938.040 1496.000 939.440 ;
        RECT 4.000 935.360 1496.000 938.040 ;
        RECT 4.000 933.960 1495.600 935.360 ;
        RECT 4.000 925.160 1496.000 933.960 ;
        RECT 4.400 923.760 1496.000 925.160 ;
        RECT 4.000 914.960 1496.000 923.760 ;
        RECT 4.000 913.560 1495.600 914.960 ;
        RECT 4.000 910.200 1496.000 913.560 ;
        RECT 4.400 908.800 1496.000 910.200 ;
        RECT 4.000 895.920 1496.000 908.800 ;
        RECT 4.400 894.560 1496.000 895.920 ;
        RECT 4.400 894.520 1495.600 894.560 ;
        RECT 4.000 893.160 1495.600 894.520 ;
        RECT 4.000 881.640 1496.000 893.160 ;
        RECT 4.400 880.240 1496.000 881.640 ;
        RECT 4.000 874.160 1496.000 880.240 ;
        RECT 4.000 872.760 1495.600 874.160 ;
        RECT 4.000 866.680 1496.000 872.760 ;
        RECT 4.400 865.280 1496.000 866.680 ;
        RECT 4.000 853.080 1496.000 865.280 ;
        RECT 4.000 852.400 1495.600 853.080 ;
        RECT 4.400 851.680 1495.600 852.400 ;
        RECT 4.400 851.000 1496.000 851.680 ;
        RECT 4.000 837.440 1496.000 851.000 ;
        RECT 4.400 836.040 1496.000 837.440 ;
        RECT 4.000 832.680 1496.000 836.040 ;
        RECT 4.000 831.280 1495.600 832.680 ;
        RECT 4.000 823.160 1496.000 831.280 ;
        RECT 4.400 821.760 1496.000 823.160 ;
        RECT 4.000 812.280 1496.000 821.760 ;
        RECT 4.000 810.880 1495.600 812.280 ;
        RECT 4.000 808.200 1496.000 810.880 ;
        RECT 4.400 806.800 1496.000 808.200 ;
        RECT 4.000 793.920 1496.000 806.800 ;
        RECT 4.400 792.520 1496.000 793.920 ;
        RECT 4.000 791.880 1496.000 792.520 ;
        RECT 4.000 790.480 1495.600 791.880 ;
        RECT 4.000 779.640 1496.000 790.480 ;
        RECT 4.400 778.240 1496.000 779.640 ;
        RECT 4.000 771.480 1496.000 778.240 ;
        RECT 4.000 770.080 1495.600 771.480 ;
        RECT 4.000 764.680 1496.000 770.080 ;
        RECT 4.400 763.280 1496.000 764.680 ;
        RECT 4.000 750.400 1496.000 763.280 ;
        RECT 4.400 749.000 1495.600 750.400 ;
        RECT 4.000 735.440 1496.000 749.000 ;
        RECT 4.400 734.040 1496.000 735.440 ;
        RECT 4.000 730.000 1496.000 734.040 ;
        RECT 4.000 728.600 1495.600 730.000 ;
        RECT 4.000 721.160 1496.000 728.600 ;
        RECT 4.400 719.760 1496.000 721.160 ;
        RECT 4.000 709.600 1496.000 719.760 ;
        RECT 4.000 708.200 1495.600 709.600 ;
        RECT 4.000 706.880 1496.000 708.200 ;
        RECT 4.400 705.480 1496.000 706.880 ;
        RECT 4.000 691.920 1496.000 705.480 ;
        RECT 4.400 690.520 1496.000 691.920 ;
        RECT 4.000 689.200 1496.000 690.520 ;
        RECT 4.000 687.800 1495.600 689.200 ;
        RECT 4.000 677.640 1496.000 687.800 ;
        RECT 4.400 676.240 1496.000 677.640 ;
        RECT 4.000 668.800 1496.000 676.240 ;
        RECT 4.000 667.400 1495.600 668.800 ;
        RECT 4.000 662.680 1496.000 667.400 ;
        RECT 4.400 661.280 1496.000 662.680 ;
        RECT 4.000 648.400 1496.000 661.280 ;
        RECT 4.400 647.720 1496.000 648.400 ;
        RECT 4.400 647.000 1495.600 647.720 ;
        RECT 4.000 646.320 1495.600 647.000 ;
        RECT 4.000 633.440 1496.000 646.320 ;
        RECT 4.400 632.040 1496.000 633.440 ;
        RECT 4.000 627.320 1496.000 632.040 ;
        RECT 4.000 625.920 1495.600 627.320 ;
        RECT 4.000 619.160 1496.000 625.920 ;
        RECT 4.400 617.760 1496.000 619.160 ;
        RECT 4.000 606.920 1496.000 617.760 ;
        RECT 4.000 605.520 1495.600 606.920 ;
        RECT 4.000 604.880 1496.000 605.520 ;
        RECT 4.400 603.480 1496.000 604.880 ;
        RECT 4.000 589.920 1496.000 603.480 ;
        RECT 4.400 588.520 1496.000 589.920 ;
        RECT 4.000 586.520 1496.000 588.520 ;
        RECT 4.000 585.120 1495.600 586.520 ;
        RECT 4.000 575.640 1496.000 585.120 ;
        RECT 4.400 574.240 1496.000 575.640 ;
        RECT 4.000 565.440 1496.000 574.240 ;
        RECT 4.000 564.040 1495.600 565.440 ;
        RECT 4.000 560.680 1496.000 564.040 ;
        RECT 4.400 559.280 1496.000 560.680 ;
        RECT 4.000 546.400 1496.000 559.280 ;
        RECT 4.400 545.040 1496.000 546.400 ;
        RECT 4.400 545.000 1495.600 545.040 ;
        RECT 4.000 543.640 1495.600 545.000 ;
        RECT 4.000 532.120 1496.000 543.640 ;
        RECT 4.400 530.720 1496.000 532.120 ;
        RECT 4.000 524.640 1496.000 530.720 ;
        RECT 4.000 523.240 1495.600 524.640 ;
        RECT 4.000 517.160 1496.000 523.240 ;
        RECT 4.400 515.760 1496.000 517.160 ;
        RECT 4.000 504.240 1496.000 515.760 ;
        RECT 4.000 502.880 1495.600 504.240 ;
        RECT 4.400 502.840 1495.600 502.880 ;
        RECT 4.400 501.480 1496.000 502.840 ;
        RECT 4.000 487.920 1496.000 501.480 ;
        RECT 4.400 486.520 1496.000 487.920 ;
        RECT 4.000 483.840 1496.000 486.520 ;
        RECT 4.000 482.440 1495.600 483.840 ;
        RECT 4.000 473.640 1496.000 482.440 ;
        RECT 4.400 472.240 1496.000 473.640 ;
        RECT 4.000 462.760 1496.000 472.240 ;
        RECT 4.000 461.360 1495.600 462.760 ;
        RECT 4.000 458.680 1496.000 461.360 ;
        RECT 4.400 457.280 1496.000 458.680 ;
        RECT 4.000 444.400 1496.000 457.280 ;
        RECT 4.400 443.000 1496.000 444.400 ;
        RECT 4.000 442.360 1496.000 443.000 ;
        RECT 4.000 440.960 1495.600 442.360 ;
        RECT 4.000 430.120 1496.000 440.960 ;
        RECT 4.400 428.720 1496.000 430.120 ;
        RECT 4.000 421.960 1496.000 428.720 ;
        RECT 4.000 420.560 1495.600 421.960 ;
        RECT 4.000 415.160 1496.000 420.560 ;
        RECT 4.400 413.760 1496.000 415.160 ;
        RECT 4.000 401.560 1496.000 413.760 ;
        RECT 4.000 400.880 1495.600 401.560 ;
        RECT 4.400 400.160 1495.600 400.880 ;
        RECT 4.400 399.480 1496.000 400.160 ;
        RECT 4.000 385.920 1496.000 399.480 ;
        RECT 4.400 384.520 1496.000 385.920 ;
        RECT 4.000 380.480 1496.000 384.520 ;
        RECT 4.000 379.080 1495.600 380.480 ;
        RECT 4.000 371.640 1496.000 379.080 ;
        RECT 4.400 370.240 1496.000 371.640 ;
        RECT 4.000 360.080 1496.000 370.240 ;
        RECT 4.000 358.680 1495.600 360.080 ;
        RECT 4.000 357.360 1496.000 358.680 ;
        RECT 4.400 355.960 1496.000 357.360 ;
        RECT 4.000 342.400 1496.000 355.960 ;
        RECT 4.400 341.000 1496.000 342.400 ;
        RECT 4.000 339.680 1496.000 341.000 ;
        RECT 4.000 338.280 1495.600 339.680 ;
        RECT 4.000 328.120 1496.000 338.280 ;
        RECT 4.400 326.720 1496.000 328.120 ;
        RECT 4.000 319.280 1496.000 326.720 ;
        RECT 4.000 317.880 1495.600 319.280 ;
        RECT 4.000 313.160 1496.000 317.880 ;
        RECT 4.400 311.760 1496.000 313.160 ;
        RECT 4.000 298.880 1496.000 311.760 ;
        RECT 4.400 297.480 1495.600 298.880 ;
        RECT 4.000 283.920 1496.000 297.480 ;
        RECT 4.400 282.520 1496.000 283.920 ;
        RECT 4.000 277.800 1496.000 282.520 ;
        RECT 4.000 276.400 1495.600 277.800 ;
        RECT 4.000 269.640 1496.000 276.400 ;
        RECT 4.400 268.240 1496.000 269.640 ;
        RECT 4.000 257.400 1496.000 268.240 ;
        RECT 4.000 256.000 1495.600 257.400 ;
        RECT 4.000 255.360 1496.000 256.000 ;
        RECT 4.400 253.960 1496.000 255.360 ;
        RECT 4.000 240.400 1496.000 253.960 ;
        RECT 4.400 239.000 1496.000 240.400 ;
        RECT 4.000 237.000 1496.000 239.000 ;
        RECT 4.000 235.600 1495.600 237.000 ;
        RECT 4.000 226.120 1496.000 235.600 ;
        RECT 4.400 224.720 1496.000 226.120 ;
        RECT 4.000 216.600 1496.000 224.720 ;
        RECT 4.000 215.200 1495.600 216.600 ;
        RECT 4.000 211.160 1496.000 215.200 ;
        RECT 4.400 209.760 1496.000 211.160 ;
        RECT 4.000 196.880 1496.000 209.760 ;
        RECT 4.400 195.520 1496.000 196.880 ;
        RECT 4.400 195.480 1495.600 195.520 ;
        RECT 4.000 194.120 1495.600 195.480 ;
        RECT 4.000 182.600 1496.000 194.120 ;
        RECT 4.400 181.200 1496.000 182.600 ;
        RECT 4.000 175.120 1496.000 181.200 ;
        RECT 4.000 173.720 1495.600 175.120 ;
        RECT 4.000 167.640 1496.000 173.720 ;
        RECT 4.400 166.240 1496.000 167.640 ;
        RECT 4.000 154.720 1496.000 166.240 ;
        RECT 4.000 153.360 1495.600 154.720 ;
        RECT 4.400 153.320 1495.600 153.360 ;
        RECT 4.400 151.960 1496.000 153.320 ;
        RECT 4.000 138.400 1496.000 151.960 ;
        RECT 4.400 137.000 1496.000 138.400 ;
        RECT 4.000 134.320 1496.000 137.000 ;
        RECT 4.000 132.920 1495.600 134.320 ;
        RECT 4.000 124.120 1496.000 132.920 ;
        RECT 4.400 122.720 1496.000 124.120 ;
        RECT 4.000 113.920 1496.000 122.720 ;
        RECT 4.000 112.520 1495.600 113.920 ;
        RECT 4.000 109.160 1496.000 112.520 ;
        RECT 4.400 107.760 1496.000 109.160 ;
        RECT 4.000 94.880 1496.000 107.760 ;
        RECT 4.400 93.480 1496.000 94.880 ;
        RECT 4.000 92.840 1496.000 93.480 ;
        RECT 4.000 91.440 1495.600 92.840 ;
        RECT 4.000 80.600 1496.000 91.440 ;
        RECT 4.400 79.200 1496.000 80.600 ;
        RECT 4.000 72.440 1496.000 79.200 ;
        RECT 4.000 71.040 1495.600 72.440 ;
        RECT 4.000 65.640 1496.000 71.040 ;
        RECT 4.400 64.240 1496.000 65.640 ;
        RECT 4.000 52.040 1496.000 64.240 ;
        RECT 4.000 51.360 1495.600 52.040 ;
        RECT 4.400 50.640 1495.600 51.360 ;
        RECT 4.400 49.960 1496.000 50.640 ;
        RECT 4.000 36.400 1496.000 49.960 ;
        RECT 4.400 35.000 1496.000 36.400 ;
        RECT 4.000 31.640 1496.000 35.000 ;
        RECT 4.000 30.240 1495.600 31.640 ;
        RECT 4.000 22.120 1496.000 30.240 ;
        RECT 4.400 20.720 1496.000 22.120 ;
        RECT 4.000 11.240 1496.000 20.720 ;
        RECT 4.000 9.840 1495.600 11.240 ;
        RECT 4.000 7.840 1496.000 9.840 ;
        RECT 4.400 6.975 1496.000 7.840 ;
      LAYER met4 ;
        RECT 212.815 10.240 251.040 1486.305 ;
        RECT 253.440 10.240 327.840 1486.305 ;
        RECT 330.240 10.240 404.640 1486.305 ;
        RECT 407.040 10.240 481.440 1486.305 ;
        RECT 483.840 10.240 558.240 1486.305 ;
        RECT 560.640 10.240 635.040 1486.305 ;
        RECT 637.440 10.240 711.840 1486.305 ;
        RECT 714.240 10.240 788.640 1486.305 ;
        RECT 791.040 10.240 865.440 1486.305 ;
        RECT 867.840 10.240 942.240 1486.305 ;
        RECT 944.640 10.240 1019.040 1486.305 ;
        RECT 1021.440 10.240 1068.745 1486.305 ;
        RECT 212.815 9.695 1068.745 10.240 ;
  END
END core
END LIBRARY

