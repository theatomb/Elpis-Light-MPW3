VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 1496.000 8.190 1500.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 8.880 1500.000 9.480 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.510 1496.000 1346.790 1500.000 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 0.000 1233.630 4.000 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.960 4.000 1271.560 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1252.600 1500.000 1253.200 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1270.960 1500.000 1271.560 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.110 0.000 1282.390 4.000 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 0.000 1298.490 4.000 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1325.360 4.000 1325.960 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 0.000 1314.590 4.000 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.510 0.000 1346.790 4.000 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.610 0.000 1362.890 4.000 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 0.000 1378.990 4.000 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1362.080 4.000 1362.680 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1325.360 1500.000 1325.960 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1398.800 4.000 1399.400 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 1496.000 1411.190 1500.000 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1417.160 4.000 1417.760 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1453.880 4.000 1454.480 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 0.000 1427.290 4.000 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1343.720 1500.000 1344.320 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.110 1496.000 1443.390 1500.000 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.210 1496.000 1459.490 1500.000 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1398.800 1500.000 1399.400 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.210 0.000 1459.490 4.000 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1435.520 1500.000 1436.120 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 0.000 1475.590 4.000 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1490.600 4.000 1491.200 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1490.600 1500.000 1491.200 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 338.000 1500.000 338.600 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 1496.000 427.250 1500.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 392.400 1500.000 393.000 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 1496.000 491.650 1500.000 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 484.200 1500.000 484.800 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 26.560 1500.000 27.160 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 502.560 1500.000 503.160 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 1496.000 588.710 1500.000 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 575.320 1500.000 575.920 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 612.040 1500.000 612.640 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 1496.000 669.210 1500.000 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 630.400 1500.000 631.000 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 1496.000 733.610 1500.000 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 1496.000 201.390 1500.000 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 1496.000 766.270 1500.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 1496.000 782.370 1500.000 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 703.840 1500.000 704.440 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 1496.000 798.470 1500.000 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 0.000 556.510 4.000 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 1496.000 814.570 1500.000 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 776.600 1500.000 777.200 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 63.280 1500.000 63.880 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 740.560 4.000 741.160 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 4.000 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 1496.000 878.970 1500.000 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 831.680 1500.000 832.280 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 0.000 685.310 4.000 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 868.400 1500.000 869.000 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 0.000 701.410 4.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 81.640 1500.000 82.240 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 1496.000 943.370 1500.000 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 905.120 1500.000 905.720 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 1496.000 959.470 1500.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 923.480 1500.000 924.080 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.680 4.000 832.280 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.760 4.000 887.360 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 959.520 1500.000 960.120 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 1496.000 266.250 1500.000 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 923.480 4.000 924.080 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 959.520 4.000 960.120 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 0.000 830.670 4.000 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 977.880 1500.000 978.480 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 0.000 846.770 4.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 996.240 1500.000 996.840 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.960 4.000 1033.560 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1051.320 4.000 1051.920 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1069.680 4.000 1070.280 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 0.000 927.270 4.000 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 0.000 959.470 4.000 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 0.000 975.570 4.000 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 1496.000 1088.730 1500.000 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 0.000 1024.330 4.000 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1051.320 1500.000 1051.920 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1088.040 1500.000 1088.640 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 118.360 1500.000 118.960 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1106.400 4.000 1107.000 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 1496.000 1120.930 1500.000 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1124.760 1500.000 1125.360 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 0.000 1104.830 4.000 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 1496.000 1153.130 1500.000 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.760 4.000 1125.360 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 1496.000 1185.330 1500.000 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 1496.000 1201.430 1500.000 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 1496.000 1249.730 1500.000 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.160 4.000 1179.760 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 1496.000 1266.290 1500.000 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.110 1496.000 1282.390 1500.000 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 0.000 1217.530 4.000 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1215.880 1500.000 1216.480 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 1496.000 1330.690 1500.000 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 246.200 1500.000 246.800 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 282.920 1500.000 283.520 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 356.360 1500.000 356.960 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 1496.000 443.350 1500.000 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 447.480 1500.000 448.080 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 1496.000 524.310 1500.000 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 520.920 1500.000 521.520 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1496.000 604.810 1500.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 593.680 1500.000 594.280 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 1496.000 620.910 1500.000 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 1496.000 685.310 1500.000 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 648.760 1500.000 649.360 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 44.920 1500.000 45.520 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 667.120 1500.000 667.720 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 100.000 1500.000 100.600 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 136.720 1500.000 137.320 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 1496.000 314.550 1500.000 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 173.440 1500.000 174.040 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 1496.000 72.590 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 1496.000 104.790 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 1496.000 120.890 1500.000 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 1496.000 88.690 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 1496.000 136.990 1500.000 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 264.560 1500.000 265.160 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 301.280 1500.000 301.880 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 1496.000 395.050 1500.000 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 374.720 1500.000 375.320 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 410.760 1500.000 411.360 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 1496.000 508.210 1500.000 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 1496.000 540.410 1500.000 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 1496.000 217.490 1500.000 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 1496.000 233.590 1500.000 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 155.080 1500.000 155.680 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 191.800 1500.000 192.400 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 1496.000 153.090 1500.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.240 4.000 1234.840 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1252.600 4.000 1253.200 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1289.320 4.000 1289.920 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 0.000 1249.730 4.000 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 0.000 1266.290 4.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1289.320 1500.000 1289.920 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1307.680 4.000 1308.280 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.720 4.000 1344.320 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 0.000 1330.690 4.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1307.680 1500.000 1308.280 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 1496.000 330.650 1500.000 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.610 1496.000 1362.890 1500.000 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.810 0.000 1395.090 4.000 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 1496.000 1378.990 1500.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.810 1496.000 1395.090 1500.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 1496.000 1427.290 1500.000 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1435.520 4.000 1436.120 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 0.000 1411.190 4.000 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.110 0.000 1443.390 4.000 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1362.080 1500.000 1362.680 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 1496.000 362.850 1500.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1380.440 1500.000 1381.040 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 1496.000 1475.590 1500.000 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 1496.000 1491.690 1500.000 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1417.160 1500.000 1417.760 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1453.880 1500.000 1454.480 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.240 4.000 1472.840 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1472.240 1500.000 1472.840 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 0.000 1491.690 4.000 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 1496.000 378.950 1500.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 1496.000 411.150 1500.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 1496.000 459.450 1500.000 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 429.120 1500.000 429.720 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 465.840 1500.000 466.440 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 1496.000 185.290 1500.000 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 1496.000 572.610 1500.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.280 4.000 539.880 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 1496.000 637.010 1500.000 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 1496.000 701.410 1500.000 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 722.200 1500.000 722.800 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 740.560 1500.000 741.160 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 1496.000 830.670 1500.000 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 758.920 1500.000 759.520 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 1496.000 846.770 1500.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 1496.000 862.870 1500.000 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 794.960 1500.000 795.560 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 813.320 1500.000 813.920 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 0.000 653.110 4.000 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 4.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 1496.000 895.070 1500.000 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 850.040 1500.000 850.640 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 1496.000 911.170 1500.000 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 886.760 1500.000 887.360 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 1496.000 927.270 1500.000 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 1496.000 249.690 1500.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.960 4.000 795.560 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 0.000 717.510 4.000 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 1496.000 975.570 1500.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 0.000 798.470 4.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 868.400 4.000 869.000 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 941.840 1500.000 942.440 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.120 4.000 905.720 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 1496.000 991.670 1500.000 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.880 4.000 978.480 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1496.000 1008.230 1500.000 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 1496.000 1024.330 1500.000 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1496.000 1040.430 1500.000 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 1496.000 1056.530 1500.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1014.600 4.000 1015.200 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 0.000 878.970 4.000 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 0.000 895.070 4.000 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 1496.000 282.350 1500.000 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1496.000 1072.630 1500.000 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 0.000 911.170 4.000 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 0.000 943.370 4.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1014.600 1500.000 1015.200 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 0.000 991.670 4.000 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1032.960 1500.000 1033.560 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 0.000 1040.430 4.000 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1069.680 1500.000 1070.280 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 1496.000 1104.830 1500.000 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1106.400 1500.000 1107.000 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1142.440 1500.000 1143.040 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 1496.000 1137.030 1500.000 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 1496.000 1169.230 1500.000 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1160.800 1500.000 1161.400 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1179.160 1500.000 1179.760 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1496.000 1217.530 1500.000 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1496.000 1233.630 1500.000 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1160.800 4.000 1161.400 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1197.520 4.000 1198.120 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 0.000 1169.230 4.000 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 0.000 1185.330 4.000 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1197.520 1500.000 1198.120 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 1496.000 1298.490 1500.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 1496.000 1314.590 1500.000 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1215.880 4.000 1216.480 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1234.240 1500.000 1234.840 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 209.480 1500.000 210.080 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 1496.000 40.390 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 1496.000 56.490 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 1496.000 169.190 1500.000 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 1496.000 346.750 1500.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 319.640 1500.000 320.240 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 1496.000 475.550 1500.000 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 1496.000 556.510 1500.000 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 539.280 1500.000 539.880 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 557.640 1500.000 558.240 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 1496.000 653.110 1500.000 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 4.000 594.280 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 1496.000 717.510 1500.000 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 1496.000 749.710 1500.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.120 4.000 667.720 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 685.480 1500.000 686.080 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 1496.000 298.450 1500.000 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 227.840 1500.000 228.440 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 1496.000 24.290 1500.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 7.225 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.080 1488.080 ;
      LAYER met2 ;
        RECT 6.990 1495.720 7.630 1496.410 ;
        RECT 8.470 1495.720 23.730 1496.410 ;
        RECT 24.570 1495.720 39.830 1496.410 ;
        RECT 40.670 1495.720 55.930 1496.410 ;
        RECT 56.770 1495.720 72.030 1496.410 ;
        RECT 72.870 1495.720 88.130 1496.410 ;
        RECT 88.970 1495.720 104.230 1496.410 ;
        RECT 105.070 1495.720 120.330 1496.410 ;
        RECT 121.170 1495.720 136.430 1496.410 ;
        RECT 137.270 1495.720 152.530 1496.410 ;
        RECT 153.370 1495.720 168.630 1496.410 ;
        RECT 169.470 1495.720 184.730 1496.410 ;
        RECT 185.570 1495.720 200.830 1496.410 ;
        RECT 201.670 1495.720 216.930 1496.410 ;
        RECT 217.770 1495.720 233.030 1496.410 ;
        RECT 233.870 1495.720 249.130 1496.410 ;
        RECT 249.970 1495.720 265.690 1496.410 ;
        RECT 266.530 1495.720 281.790 1496.410 ;
        RECT 282.630 1495.720 297.890 1496.410 ;
        RECT 298.730 1495.720 313.990 1496.410 ;
        RECT 314.830 1495.720 330.090 1496.410 ;
        RECT 330.930 1495.720 346.190 1496.410 ;
        RECT 347.030 1495.720 362.290 1496.410 ;
        RECT 363.130 1495.720 378.390 1496.410 ;
        RECT 379.230 1495.720 394.490 1496.410 ;
        RECT 395.330 1495.720 410.590 1496.410 ;
        RECT 411.430 1495.720 426.690 1496.410 ;
        RECT 427.530 1495.720 442.790 1496.410 ;
        RECT 443.630 1495.720 458.890 1496.410 ;
        RECT 459.730 1495.720 474.990 1496.410 ;
        RECT 475.830 1495.720 491.090 1496.410 ;
        RECT 491.930 1495.720 507.650 1496.410 ;
        RECT 508.490 1495.720 523.750 1496.410 ;
        RECT 524.590 1495.720 539.850 1496.410 ;
        RECT 540.690 1495.720 555.950 1496.410 ;
        RECT 556.790 1495.720 572.050 1496.410 ;
        RECT 572.890 1495.720 588.150 1496.410 ;
        RECT 588.990 1495.720 604.250 1496.410 ;
        RECT 605.090 1495.720 620.350 1496.410 ;
        RECT 621.190 1495.720 636.450 1496.410 ;
        RECT 637.290 1495.720 652.550 1496.410 ;
        RECT 653.390 1495.720 668.650 1496.410 ;
        RECT 669.490 1495.720 684.750 1496.410 ;
        RECT 685.590 1495.720 700.850 1496.410 ;
        RECT 701.690 1495.720 716.950 1496.410 ;
        RECT 717.790 1495.720 733.050 1496.410 ;
        RECT 733.890 1495.720 749.150 1496.410 ;
        RECT 749.990 1495.720 765.710 1496.410 ;
        RECT 766.550 1495.720 781.810 1496.410 ;
        RECT 782.650 1495.720 797.910 1496.410 ;
        RECT 798.750 1495.720 814.010 1496.410 ;
        RECT 814.850 1495.720 830.110 1496.410 ;
        RECT 830.950 1495.720 846.210 1496.410 ;
        RECT 847.050 1495.720 862.310 1496.410 ;
        RECT 863.150 1495.720 878.410 1496.410 ;
        RECT 879.250 1495.720 894.510 1496.410 ;
        RECT 895.350 1495.720 910.610 1496.410 ;
        RECT 911.450 1495.720 926.710 1496.410 ;
        RECT 927.550 1495.720 942.810 1496.410 ;
        RECT 943.650 1495.720 958.910 1496.410 ;
        RECT 959.750 1495.720 975.010 1496.410 ;
        RECT 975.850 1495.720 991.110 1496.410 ;
        RECT 991.950 1495.720 1007.670 1496.410 ;
        RECT 1008.510 1495.720 1023.770 1496.410 ;
        RECT 1024.610 1495.720 1039.870 1496.410 ;
        RECT 1040.710 1495.720 1055.970 1496.410 ;
        RECT 1056.810 1495.720 1072.070 1496.410 ;
        RECT 1072.910 1495.720 1088.170 1496.410 ;
        RECT 1089.010 1495.720 1104.270 1496.410 ;
        RECT 1105.110 1495.720 1120.370 1496.410 ;
        RECT 1121.210 1495.720 1136.470 1496.410 ;
        RECT 1137.310 1495.720 1152.570 1496.410 ;
        RECT 1153.410 1495.720 1168.670 1496.410 ;
        RECT 1169.510 1495.720 1184.770 1496.410 ;
        RECT 1185.610 1495.720 1200.870 1496.410 ;
        RECT 1201.710 1495.720 1216.970 1496.410 ;
        RECT 1217.810 1495.720 1233.070 1496.410 ;
        RECT 1233.910 1495.720 1249.170 1496.410 ;
        RECT 1250.010 1495.720 1265.730 1496.410 ;
        RECT 1266.570 1495.720 1281.830 1496.410 ;
        RECT 1282.670 1495.720 1297.930 1496.410 ;
        RECT 1298.770 1495.720 1314.030 1496.410 ;
        RECT 1314.870 1495.720 1330.130 1496.410 ;
        RECT 1330.970 1495.720 1346.230 1496.410 ;
        RECT 1347.070 1495.720 1362.330 1496.410 ;
        RECT 1363.170 1495.720 1378.430 1496.410 ;
        RECT 1379.270 1495.720 1394.530 1496.410 ;
        RECT 1395.370 1495.720 1410.630 1496.410 ;
        RECT 1411.470 1495.720 1426.730 1496.410 ;
        RECT 1427.570 1495.720 1442.830 1496.410 ;
        RECT 1443.670 1495.720 1458.930 1496.410 ;
        RECT 1459.770 1495.720 1475.030 1496.410 ;
        RECT 1475.870 1495.720 1491.130 1496.410 ;
        RECT 6.990 4.280 1491.680 1495.720 ;
        RECT 6.990 3.670 7.630 4.280 ;
        RECT 8.470 3.670 23.730 4.280 ;
        RECT 24.570 3.670 39.830 4.280 ;
        RECT 40.670 3.670 55.930 4.280 ;
        RECT 56.770 3.670 72.030 4.280 ;
        RECT 72.870 3.670 88.130 4.280 ;
        RECT 88.970 3.670 104.230 4.280 ;
        RECT 105.070 3.670 120.330 4.280 ;
        RECT 121.170 3.670 136.430 4.280 ;
        RECT 137.270 3.670 152.530 4.280 ;
        RECT 153.370 3.670 168.630 4.280 ;
        RECT 169.470 3.670 184.730 4.280 ;
        RECT 185.570 3.670 200.830 4.280 ;
        RECT 201.670 3.670 216.930 4.280 ;
        RECT 217.770 3.670 233.030 4.280 ;
        RECT 233.870 3.670 249.130 4.280 ;
        RECT 249.970 3.670 265.690 4.280 ;
        RECT 266.530 3.670 281.790 4.280 ;
        RECT 282.630 3.670 297.890 4.280 ;
        RECT 298.730 3.670 313.990 4.280 ;
        RECT 314.830 3.670 330.090 4.280 ;
        RECT 330.930 3.670 346.190 4.280 ;
        RECT 347.030 3.670 362.290 4.280 ;
        RECT 363.130 3.670 378.390 4.280 ;
        RECT 379.230 3.670 394.490 4.280 ;
        RECT 395.330 3.670 410.590 4.280 ;
        RECT 411.430 3.670 426.690 4.280 ;
        RECT 427.530 3.670 442.790 4.280 ;
        RECT 443.630 3.670 458.890 4.280 ;
        RECT 459.730 3.670 474.990 4.280 ;
        RECT 475.830 3.670 491.090 4.280 ;
        RECT 491.930 3.670 507.650 4.280 ;
        RECT 508.490 3.670 523.750 4.280 ;
        RECT 524.590 3.670 539.850 4.280 ;
        RECT 540.690 3.670 555.950 4.280 ;
        RECT 556.790 3.670 572.050 4.280 ;
        RECT 572.890 3.670 588.150 4.280 ;
        RECT 588.990 3.670 604.250 4.280 ;
        RECT 605.090 3.670 620.350 4.280 ;
        RECT 621.190 3.670 636.450 4.280 ;
        RECT 637.290 3.670 652.550 4.280 ;
        RECT 653.390 3.670 668.650 4.280 ;
        RECT 669.490 3.670 684.750 4.280 ;
        RECT 685.590 3.670 700.850 4.280 ;
        RECT 701.690 3.670 716.950 4.280 ;
        RECT 717.790 3.670 733.050 4.280 ;
        RECT 733.890 3.670 749.150 4.280 ;
        RECT 749.990 3.670 765.710 4.280 ;
        RECT 766.550 3.670 781.810 4.280 ;
        RECT 782.650 3.670 797.910 4.280 ;
        RECT 798.750 3.670 814.010 4.280 ;
        RECT 814.850 3.670 830.110 4.280 ;
        RECT 830.950 3.670 846.210 4.280 ;
        RECT 847.050 3.670 862.310 4.280 ;
        RECT 863.150 3.670 878.410 4.280 ;
        RECT 879.250 3.670 894.510 4.280 ;
        RECT 895.350 3.670 910.610 4.280 ;
        RECT 911.450 3.670 926.710 4.280 ;
        RECT 927.550 3.670 942.810 4.280 ;
        RECT 943.650 3.670 958.910 4.280 ;
        RECT 959.750 3.670 975.010 4.280 ;
        RECT 975.850 3.670 991.110 4.280 ;
        RECT 991.950 3.670 1007.670 4.280 ;
        RECT 1008.510 3.670 1023.770 4.280 ;
        RECT 1024.610 3.670 1039.870 4.280 ;
        RECT 1040.710 3.670 1055.970 4.280 ;
        RECT 1056.810 3.670 1072.070 4.280 ;
        RECT 1072.910 3.670 1088.170 4.280 ;
        RECT 1089.010 3.670 1104.270 4.280 ;
        RECT 1105.110 3.670 1120.370 4.280 ;
        RECT 1121.210 3.670 1136.470 4.280 ;
        RECT 1137.310 3.670 1152.570 4.280 ;
        RECT 1153.410 3.670 1168.670 4.280 ;
        RECT 1169.510 3.670 1184.770 4.280 ;
        RECT 1185.610 3.670 1200.870 4.280 ;
        RECT 1201.710 3.670 1216.970 4.280 ;
        RECT 1217.810 3.670 1233.070 4.280 ;
        RECT 1233.910 3.670 1249.170 4.280 ;
        RECT 1250.010 3.670 1265.730 4.280 ;
        RECT 1266.570 3.670 1281.830 4.280 ;
        RECT 1282.670 3.670 1297.930 4.280 ;
        RECT 1298.770 3.670 1314.030 4.280 ;
        RECT 1314.870 3.670 1330.130 4.280 ;
        RECT 1330.970 3.670 1346.230 4.280 ;
        RECT 1347.070 3.670 1362.330 4.280 ;
        RECT 1363.170 3.670 1378.430 4.280 ;
        RECT 1379.270 3.670 1394.530 4.280 ;
        RECT 1395.370 3.670 1410.630 4.280 ;
        RECT 1411.470 3.670 1426.730 4.280 ;
        RECT 1427.570 3.670 1442.830 4.280 ;
        RECT 1443.670 3.670 1458.930 4.280 ;
        RECT 1459.770 3.670 1475.030 4.280 ;
        RECT 1475.870 3.670 1491.130 4.280 ;
      LAYER met3 ;
        RECT 4.400 1490.200 1495.600 1491.065 ;
        RECT 4.000 1473.240 1496.000 1490.200 ;
        RECT 4.400 1471.840 1495.600 1473.240 ;
        RECT 4.000 1454.880 1496.000 1471.840 ;
        RECT 4.400 1453.480 1495.600 1454.880 ;
        RECT 4.000 1436.520 1496.000 1453.480 ;
        RECT 4.400 1435.120 1495.600 1436.520 ;
        RECT 4.000 1418.160 1496.000 1435.120 ;
        RECT 4.400 1416.760 1495.600 1418.160 ;
        RECT 4.000 1399.800 1496.000 1416.760 ;
        RECT 4.400 1398.400 1495.600 1399.800 ;
        RECT 4.000 1381.440 1496.000 1398.400 ;
        RECT 4.400 1380.040 1495.600 1381.440 ;
        RECT 4.000 1363.080 1496.000 1380.040 ;
        RECT 4.400 1361.680 1495.600 1363.080 ;
        RECT 4.000 1344.720 1496.000 1361.680 ;
        RECT 4.400 1343.320 1495.600 1344.720 ;
        RECT 4.000 1326.360 1496.000 1343.320 ;
        RECT 4.400 1324.960 1495.600 1326.360 ;
        RECT 4.000 1308.680 1496.000 1324.960 ;
        RECT 4.400 1307.280 1495.600 1308.680 ;
        RECT 4.000 1290.320 1496.000 1307.280 ;
        RECT 4.400 1288.920 1495.600 1290.320 ;
        RECT 4.000 1271.960 1496.000 1288.920 ;
        RECT 4.400 1270.560 1495.600 1271.960 ;
        RECT 4.000 1253.600 1496.000 1270.560 ;
        RECT 4.400 1252.200 1495.600 1253.600 ;
        RECT 4.000 1235.240 1496.000 1252.200 ;
        RECT 4.400 1233.840 1495.600 1235.240 ;
        RECT 4.000 1216.880 1496.000 1233.840 ;
        RECT 4.400 1215.480 1495.600 1216.880 ;
        RECT 4.000 1198.520 1496.000 1215.480 ;
        RECT 4.400 1197.120 1495.600 1198.520 ;
        RECT 4.000 1180.160 1496.000 1197.120 ;
        RECT 4.400 1178.760 1495.600 1180.160 ;
        RECT 4.000 1161.800 1496.000 1178.760 ;
        RECT 4.400 1160.400 1495.600 1161.800 ;
        RECT 4.000 1143.440 1496.000 1160.400 ;
        RECT 4.400 1142.040 1495.600 1143.440 ;
        RECT 4.000 1125.760 1496.000 1142.040 ;
        RECT 4.400 1124.360 1495.600 1125.760 ;
        RECT 4.000 1107.400 1496.000 1124.360 ;
        RECT 4.400 1106.000 1495.600 1107.400 ;
        RECT 4.000 1089.040 1496.000 1106.000 ;
        RECT 4.400 1087.640 1495.600 1089.040 ;
        RECT 4.000 1070.680 1496.000 1087.640 ;
        RECT 4.400 1069.280 1495.600 1070.680 ;
        RECT 4.000 1052.320 1496.000 1069.280 ;
        RECT 4.400 1050.920 1495.600 1052.320 ;
        RECT 4.000 1033.960 1496.000 1050.920 ;
        RECT 4.400 1032.560 1495.600 1033.960 ;
        RECT 4.000 1015.600 1496.000 1032.560 ;
        RECT 4.400 1014.200 1495.600 1015.600 ;
        RECT 4.000 997.240 1496.000 1014.200 ;
        RECT 4.400 995.840 1495.600 997.240 ;
        RECT 4.000 978.880 1496.000 995.840 ;
        RECT 4.400 977.480 1495.600 978.880 ;
        RECT 4.000 960.520 1496.000 977.480 ;
        RECT 4.400 959.120 1495.600 960.520 ;
        RECT 4.000 942.840 1496.000 959.120 ;
        RECT 4.400 941.440 1495.600 942.840 ;
        RECT 4.000 924.480 1496.000 941.440 ;
        RECT 4.400 923.080 1495.600 924.480 ;
        RECT 4.000 906.120 1496.000 923.080 ;
        RECT 4.400 904.720 1495.600 906.120 ;
        RECT 4.000 887.760 1496.000 904.720 ;
        RECT 4.400 886.360 1495.600 887.760 ;
        RECT 4.000 869.400 1496.000 886.360 ;
        RECT 4.400 868.000 1495.600 869.400 ;
        RECT 4.000 851.040 1496.000 868.000 ;
        RECT 4.400 849.640 1495.600 851.040 ;
        RECT 4.000 832.680 1496.000 849.640 ;
        RECT 4.400 831.280 1495.600 832.680 ;
        RECT 4.000 814.320 1496.000 831.280 ;
        RECT 4.400 812.920 1495.600 814.320 ;
        RECT 4.000 795.960 1496.000 812.920 ;
        RECT 4.400 794.560 1495.600 795.960 ;
        RECT 4.000 777.600 1496.000 794.560 ;
        RECT 4.400 776.200 1495.600 777.600 ;
        RECT 4.000 759.920 1496.000 776.200 ;
        RECT 4.400 758.520 1495.600 759.920 ;
        RECT 4.000 741.560 1496.000 758.520 ;
        RECT 4.400 740.160 1495.600 741.560 ;
        RECT 4.000 723.200 1496.000 740.160 ;
        RECT 4.400 721.800 1495.600 723.200 ;
        RECT 4.000 704.840 1496.000 721.800 ;
        RECT 4.400 703.440 1495.600 704.840 ;
        RECT 4.000 686.480 1496.000 703.440 ;
        RECT 4.400 685.080 1495.600 686.480 ;
        RECT 4.000 668.120 1496.000 685.080 ;
        RECT 4.400 666.720 1495.600 668.120 ;
        RECT 4.000 649.760 1496.000 666.720 ;
        RECT 4.400 648.360 1495.600 649.760 ;
        RECT 4.000 631.400 1496.000 648.360 ;
        RECT 4.400 630.000 1495.600 631.400 ;
        RECT 4.000 613.040 1496.000 630.000 ;
        RECT 4.400 611.640 1495.600 613.040 ;
        RECT 4.000 594.680 1496.000 611.640 ;
        RECT 4.400 593.280 1495.600 594.680 ;
        RECT 4.000 576.320 1496.000 593.280 ;
        RECT 4.400 574.920 1495.600 576.320 ;
        RECT 4.000 558.640 1496.000 574.920 ;
        RECT 4.400 557.240 1495.600 558.640 ;
        RECT 4.000 540.280 1496.000 557.240 ;
        RECT 4.400 538.880 1495.600 540.280 ;
        RECT 4.000 521.920 1496.000 538.880 ;
        RECT 4.400 520.520 1495.600 521.920 ;
        RECT 4.000 503.560 1496.000 520.520 ;
        RECT 4.400 502.160 1495.600 503.560 ;
        RECT 4.000 485.200 1496.000 502.160 ;
        RECT 4.400 483.800 1495.600 485.200 ;
        RECT 4.000 466.840 1496.000 483.800 ;
        RECT 4.400 465.440 1495.600 466.840 ;
        RECT 4.000 448.480 1496.000 465.440 ;
        RECT 4.400 447.080 1495.600 448.480 ;
        RECT 4.000 430.120 1496.000 447.080 ;
        RECT 4.400 428.720 1495.600 430.120 ;
        RECT 4.000 411.760 1496.000 428.720 ;
        RECT 4.400 410.360 1495.600 411.760 ;
        RECT 4.000 393.400 1496.000 410.360 ;
        RECT 4.400 392.000 1495.600 393.400 ;
        RECT 4.000 375.720 1496.000 392.000 ;
        RECT 4.400 374.320 1495.600 375.720 ;
        RECT 4.000 357.360 1496.000 374.320 ;
        RECT 4.400 355.960 1495.600 357.360 ;
        RECT 4.000 339.000 1496.000 355.960 ;
        RECT 4.400 337.600 1495.600 339.000 ;
        RECT 4.000 320.640 1496.000 337.600 ;
        RECT 4.400 319.240 1495.600 320.640 ;
        RECT 4.000 302.280 1496.000 319.240 ;
        RECT 4.400 300.880 1495.600 302.280 ;
        RECT 4.000 283.920 1496.000 300.880 ;
        RECT 4.400 282.520 1495.600 283.920 ;
        RECT 4.000 265.560 1496.000 282.520 ;
        RECT 4.400 264.160 1495.600 265.560 ;
        RECT 4.000 247.200 1496.000 264.160 ;
        RECT 4.400 245.800 1495.600 247.200 ;
        RECT 4.000 228.840 1496.000 245.800 ;
        RECT 4.400 227.440 1495.600 228.840 ;
        RECT 4.000 210.480 1496.000 227.440 ;
        RECT 4.400 209.080 1495.600 210.480 ;
        RECT 4.000 192.800 1496.000 209.080 ;
        RECT 4.400 191.400 1495.600 192.800 ;
        RECT 4.000 174.440 1496.000 191.400 ;
        RECT 4.400 173.040 1495.600 174.440 ;
        RECT 4.000 156.080 1496.000 173.040 ;
        RECT 4.400 154.680 1495.600 156.080 ;
        RECT 4.000 137.720 1496.000 154.680 ;
        RECT 4.400 136.320 1495.600 137.720 ;
        RECT 4.000 119.360 1496.000 136.320 ;
        RECT 4.400 117.960 1495.600 119.360 ;
        RECT 4.000 101.000 1496.000 117.960 ;
        RECT 4.400 99.600 1495.600 101.000 ;
        RECT 4.000 82.640 1496.000 99.600 ;
        RECT 4.400 81.240 1495.600 82.640 ;
        RECT 4.000 64.280 1496.000 81.240 ;
        RECT 4.400 62.880 1495.600 64.280 ;
        RECT 4.000 45.920 1496.000 62.880 ;
        RECT 4.400 44.520 1495.600 45.920 ;
        RECT 4.000 27.560 1496.000 44.520 ;
        RECT 4.400 26.160 1495.600 27.560 ;
        RECT 4.000 9.880 1496.000 26.160 ;
        RECT 4.400 9.015 1495.600 9.880 ;
      LAYER met4 ;
        RECT 366.455 12.415 404.640 1485.625 ;
        RECT 407.040 12.415 481.440 1485.625 ;
        RECT 483.840 12.415 558.240 1485.625 ;
        RECT 560.640 12.415 635.040 1485.625 ;
        RECT 637.440 12.415 711.840 1485.625 ;
        RECT 714.240 12.415 788.640 1485.625 ;
        RECT 791.040 12.415 865.440 1485.625 ;
        RECT 867.840 12.415 942.240 1485.625 ;
        RECT 944.640 12.415 1019.040 1485.625 ;
        RECT 1021.440 12.415 1092.665 1485.625 ;
  END
END core
END LIBRARY

