VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_controller
  CLASS BLOCK ;
  FOREIGN chip_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN addr0_to_sram[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END addr0_to_sram[0]
  PIN addr0_to_sram[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END addr0_to_sram[10]
  PIN addr0_to_sram[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 78.240 400.000 78.840 ;
    END
  END addr0_to_sram[11]
  PIN addr0_to_sram[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END addr0_to_sram[12]
  PIN addr0_to_sram[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END addr0_to_sram[13]
  PIN addr0_to_sram[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 396.000 87.310 400.000 ;
    END
  END addr0_to_sram[14]
  PIN addr0_to_sram[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END addr0_to_sram[15]
  PIN addr0_to_sram[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 102.040 400.000 102.640 ;
    END
  END addr0_to_sram[16]
  PIN addr0_to_sram[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END addr0_to_sram[17]
  PIN addr0_to_sram[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 117.000 400.000 117.600 ;
    END
  END addr0_to_sram[18]
  PIN addr0_to_sram[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.120 400.000 123.720 ;
    END
  END addr0_to_sram[19]
  PIN addr0_to_sram[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END addr0_to_sram[1]
  PIN addr0_to_sram[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 396.000 14.630 400.000 ;
    END
  END addr0_to_sram[2]
  PIN addr0_to_sram[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END addr0_to_sram[3]
  PIN addr0_to_sram[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 26.560 400.000 27.160 ;
    END
  END addr0_to_sram[4]
  PIN addr0_to_sram[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 39.480 400.000 40.080 ;
    END
  END addr0_to_sram[5]
  PIN addr0_to_sram[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END addr0_to_sram[6]
  PIN addr0_to_sram[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 58.520 400.000 59.120 ;
    END
  END addr0_to_sram[7]
  PIN addr0_to_sram[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 63.280 400.000 63.880 ;
    END
  END addr0_to_sram[8]
  PIN addr0_to_sram[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 66.680 400.000 67.280 ;
    END
  END addr0_to_sram[9]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END addr_in[0]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END addr_in[11]
  PIN addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END addr_in[12]
  PIN addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END addr_in[13]
  PIN addr_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 92.520 400.000 93.120 ;
    END
  END addr_in[14]
  PIN addr_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END addr_in[15]
  PIN addr_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 396.000 101.110 400.000 ;
    END
  END addr_in[16]
  PIN addr_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END addr_in[17]
  PIN addr_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 396.000 118.590 400.000 ;
    END
  END addr_in[18]
  PIN addr_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END addr_in[19]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 21.120 400.000 21.720 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 27.920 400.000 28.520 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 40.840 400.000 41.440 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 396.000 47.290 400.000 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 396.000 57.870 400.000 ;
    END
  END addr_in[9]
  PIN addr_to_core_mem[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 5.480 400.000 6.080 ;
    END
  END addr_to_core_mem[0]
  PIN addr_to_core_mem[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END addr_to_core_mem[10]
  PIN addr_to_core_mem[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 79.600 400.000 80.200 ;
    END
  END addr_to_core_mem[11]
  PIN addr_to_core_mem[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 83.000 400.000 83.600 ;
    END
  END addr_to_core_mem[12]
  PIN addr_to_core_mem[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END addr_to_core_mem[13]
  PIN addr_to_core_mem[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 396.000 89.150 400.000 ;
    END
  END addr_to_core_mem[14]
  PIN addr_to_core_mem[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 97.280 400.000 97.880 ;
    END
  END addr_to_core_mem[15]
  PIN addr_to_core_mem[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END addr_to_core_mem[16]
  PIN addr_to_core_mem[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END addr_to_core_mem[17]
  PIN addr_to_core_mem[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END addr_to_core_mem[18]
  PIN addr_to_core_mem[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 125.160 400.000 125.760 ;
    END
  END addr_to_core_mem[19]
  PIN addr_to_core_mem[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END addr_to_core_mem[1]
  PIN addr_to_core_mem[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 396.000 16.010 400.000 ;
    END
  END addr_to_core_mem[2]
  PIN addr_to_core_mem[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END addr_to_core_mem[3]
  PIN addr_to_core_mem[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END addr_to_core_mem[4]
  PIN addr_to_core_mem[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 42.200 400.000 42.800 ;
    END
  END addr_to_core_mem[5]
  PIN addr_to_core_mem[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 50.360 400.000 50.960 ;
    END
  END addr_to_core_mem[6]
  PIN addr_to_core_mem[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END addr_to_core_mem[7]
  PIN addr_to_core_mem[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 396.000 49.130 400.000 ;
    END
  END addr_to_core_mem[8]
  PIN addr_to_core_mem[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.040 400.000 68.640 ;
    END
  END addr_to_core_mem[9]
  PIN clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END clk
  PIN core0_data_print[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END core0_data_print[0]
  PIN core0_data_print[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END core0_data_print[10]
  PIN core0_data_print[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 396.000 67.990 400.000 ;
    END
  END core0_data_print[11]
  PIN core0_data_print[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END core0_data_print[12]
  PIN core0_data_print[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 396.000 78.570 400.000 ;
    END
  END core0_data_print[13]
  PIN core0_data_print[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END core0_data_print[14]
  PIN core0_data_print[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 396.000 92.370 400.000 ;
    END
  END core0_data_print[15]
  PIN core0_data_print[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 104.080 400.000 104.680 ;
    END
  END core0_data_print[16]
  PIN core0_data_print[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 107.480 400.000 108.080 ;
    END
  END core0_data_print[17]
  PIN core0_data_print[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END core0_data_print[18]
  PIN core0_data_print[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END core0_data_print[19]
  PIN core0_data_print[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 8.200 400.000 8.800 ;
    END
  END core0_data_print[1]
  PIN core0_data_print[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END core0_data_print[20]
  PIN core0_data_print[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END core0_data_print[21]
  PIN core0_data_print[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END core0_data_print[22]
  PIN core0_data_print[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END core0_data_print[23]
  PIN core0_data_print[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END core0_data_print[24]
  PIN core0_data_print[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.160 400.000 159.760 ;
    END
  END core0_data_print[25]
  PIN core0_data_print[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 163.920 400.000 164.520 ;
    END
  END core0_data_print[26]
  PIN core0_data_print[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END core0_data_print[27]
  PIN core0_data_print[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END core0_data_print[28]
  PIN core0_data_print[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END core0_data_print[29]
  PIN core0_data_print[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 396.000 17.850 400.000 ;
    END
  END core0_data_print[2]
  PIN core0_data_print[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END core0_data_print[30]
  PIN core0_data_print[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 183.640 400.000 184.240 ;
    END
  END core0_data_print[31]
  PIN core0_data_print[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END core0_data_print[3]
  PIN core0_data_print[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 29.280 400.000 29.880 ;
    END
  END core0_data_print[4]
  PIN core0_data_print[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 44.240 400.000 44.840 ;
    END
  END core0_data_print[5]
  PIN core0_data_print[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END core0_data_print[6]
  PIN core0_data_print[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 396.000 40.390 400.000 ;
    END
  END core0_data_print[7]
  PIN core0_data_print[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END core0_data_print[8]
  PIN core0_data_print[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END core0_data_print[9]
  PIN csb0_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 2.080 400.000 2.680 ;
    END
  END csb0_to_sram
  PIN data_out_to_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END data_out_to_core[0]
  PIN data_out_to_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 73.480 400.000 74.080 ;
    END
  END data_out_to_core[10]
  PIN data_out_to_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END data_out_to_core[11]
  PIN data_out_to_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END data_out_to_core[12]
  PIN data_out_to_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 396.000 80.410 400.000 ;
    END
  END data_out_to_core[13]
  PIN data_out_to_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END data_out_to_core[14]
  PIN data_out_to_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 396.000 94.210 400.000 ;
    END
  END data_out_to_core[15]
  PIN data_out_to_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 396.000 102.950 400.000 ;
    END
  END data_out_to_core[16]
  PIN data_out_to_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 108.840 400.000 109.440 ;
    END
  END data_out_to_core[17]
  PIN data_out_to_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 396.000 119.970 400.000 ;
    END
  END data_out_to_core[18]
  PIN data_out_to_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END data_out_to_core[19]
  PIN data_out_to_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END data_out_to_core[1]
  PIN data_out_to_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END data_out_to_core[20]
  PIN data_out_to_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 134.680 400.000 135.280 ;
    END
  END data_out_to_core[21]
  PIN data_out_to_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 396.000 141.130 400.000 ;
    END
  END data_out_to_core[22]
  PIN data_out_to_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.840 400.000 143.440 ;
    END
  END data_out_to_core[23]
  PIN data_out_to_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END data_out_to_core[24]
  PIN data_out_to_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END data_out_to_core[25]
  PIN data_out_to_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 396.000 163.670 400.000 ;
    END
  END data_out_to_core[26]
  PIN data_out_to_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END data_out_to_core[27]
  PIN data_out_to_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 396.000 177.470 400.000 ;
    END
  END data_out_to_core[28]
  PIN data_out_to_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 176.840 400.000 177.440 ;
    END
  END data_out_to_core[29]
  PIN data_out_to_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END data_out_to_core[2]
  PIN data_out_to_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END data_out_to_core[30]
  PIN data_out_to_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END data_out_to_core[31]
  PIN data_out_to_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 23.160 400.000 23.760 ;
    END
  END data_out_to_core[3]
  PIN data_out_to_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END data_out_to_core[4]
  PIN data_out_to_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END data_out_to_core[5]
  PIN data_out_to_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 52.400 400.000 53.000 ;
    END
  END data_out_to_core[6]
  PIN data_out_to_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END data_out_to_core[7]
  PIN data_out_to_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END data_out_to_core[8]
  PIN data_out_to_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END data_out_to_core[9]
  PIN data_to_core_mem[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 6.840 400.000 7.440 ;
    END
  END data_to_core_mem[0]
  PIN data_to_core_mem[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END data_to_core_mem[10]
  PIN data_to_core_mem[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END data_to_core_mem[11]
  PIN data_to_core_mem[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END data_to_core_mem[12]
  PIN data_to_core_mem[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 396.000 82.250 400.000 ;
    END
  END data_to_core_mem[13]
  PIN data_to_core_mem[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 94.560 400.000 95.160 ;
    END
  END data_to_core_mem[14]
  PIN data_to_core_mem[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END data_to_core_mem[15]
  PIN data_to_core_mem[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END data_to_core_mem[16]
  PIN data_to_core_mem[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 396.000 111.690 400.000 ;
    END
  END data_to_core_mem[17]
  PIN data_to_core_mem[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END data_to_core_mem[18]
  PIN data_to_core_mem[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 126.520 400.000 127.120 ;
    END
  END data_to_core_mem[19]
  PIN data_to_core_mem[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 396.000 9.110 400.000 ;
    END
  END data_to_core_mem[1]
  PIN data_to_core_mem[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END data_to_core_mem[20]
  PIN data_to_core_mem[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 136.040 400.000 136.640 ;
    END
  END data_to_core_mem[21]
  PIN data_to_core_mem[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 396.000 142.510 400.000 ;
    END
  END data_to_core_mem[22]
  PIN data_to_core_mem[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 144.200 400.000 144.800 ;
    END
  END data_to_core_mem[23]
  PIN data_to_core_mem[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END data_to_core_mem[24]
  PIN data_to_core_mem[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 396.000 154.930 400.000 ;
    END
  END data_to_core_mem[25]
  PIN data_to_core_mem[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 396.000 165.050 400.000 ;
    END
  END data_to_core_mem[26]
  PIN data_to_core_mem[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END data_to_core_mem[27]
  PIN data_to_core_mem[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 175.480 400.000 176.080 ;
    END
  END data_to_core_mem[28]
  PIN data_to_core_mem[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END data_to_core_mem[29]
  PIN data_to_core_mem[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END data_to_core_mem[2]
  PIN data_to_core_mem[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END data_to_core_mem[30]
  PIN data_to_core_mem[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END data_to_core_mem[31]
  PIN data_to_core_mem[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END data_to_core_mem[3]
  PIN data_to_core_mem[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 31.320 400.000 31.920 ;
    END
  END data_to_core_mem[4]
  PIN data_to_core_mem[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 45.600 400.000 46.200 ;
    END
  END data_to_core_mem[5]
  PIN data_to_core_mem[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END data_to_core_mem[6]
  PIN data_to_core_mem[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END data_to_core_mem[7]
  PIN data_to_core_mem[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END data_to_core_mem[8]
  PIN data_to_core_mem[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END data_to_core_mem[9]
  PIN din0_to_sram[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END din0_to_sram[0]
  PIN din0_to_sram[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 396.000 62.930 400.000 ;
    END
  END din0_to_sram[10]
  PIN din0_to_sram[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END din0_to_sram[11]
  PIN din0_to_sram[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 84.360 400.000 84.960 ;
    END
  END din0_to_sram[12]
  PIN din0_to_sram[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END din0_to_sram[13]
  PIN din0_to_sram[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END din0_to_sram[14]
  PIN din0_to_sram[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END din0_to_sram[15]
  PIN din0_to_sram[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 396.000 104.330 400.000 ;
    END
  END din0_to_sram[16]
  PIN din0_to_sram[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 110.200 400.000 110.800 ;
    END
  END din0_to_sram[17]
  PIN din0_to_sram[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 396.000 121.810 400.000 ;
    END
  END din0_to_sram[18]
  PIN din0_to_sram[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 128.560 400.000 129.160 ;
    END
  END din0_to_sram[19]
  PIN din0_to_sram[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 10.240 400.000 10.840 ;
    END
  END din0_to_sram[1]
  PIN din0_to_sram[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END din0_to_sram[20]
  PIN din0_to_sram[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END din0_to_sram[21]
  PIN din0_to_sram[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END din0_to_sram[22]
  PIN din0_to_sram[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END din0_to_sram[23]
  PIN din0_to_sram[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END din0_to_sram[24]
  PIN din0_to_sram[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 396.000 156.310 400.000 ;
    END
  END din0_to_sram[25]
  PIN din0_to_sram[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END din0_to_sram[26]
  PIN din0_to_sram[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 168.680 400.000 169.280 ;
    END
  END din0_to_sram[27]
  PIN din0_to_sram[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END din0_to_sram[28]
  PIN din0_to_sram[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END din0_to_sram[29]
  PIN din0_to_sram[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 396.000 19.690 400.000 ;
    END
  END din0_to_sram[2]
  PIN din0_to_sram[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.240 400.000 180.840 ;
    END
  END din0_to_sram[30]
  PIN din0_to_sram[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END din0_to_sram[31]
  PIN din0_to_sram[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 24.520 400.000 25.120 ;
    END
  END din0_to_sram[3]
  PIN din0_to_sram[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END din0_to_sram[4]
  PIN din0_to_sram[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END din0_to_sram[5]
  PIN din0_to_sram[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 53.760 400.000 54.360 ;
    END
  END din0_to_sram[6]
  PIN din0_to_sram[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END din0_to_sram[7]
  PIN din0_to_sram[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 396.000 50.970 400.000 ;
    END
  END din0_to_sram[8]
  PIN din0_to_sram[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END din0_to_sram[9]
  PIN dout0_to_sram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END dout0_to_sram[0]
  PIN dout0_to_sram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END dout0_to_sram[10]
  PIN dout0_to_sram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 396.000 69.830 400.000 ;
    END
  END dout0_to_sram[11]
  PIN dout0_to_sram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 396.000 74.890 400.000 ;
    END
  END dout0_to_sram[12]
  PIN dout0_to_sram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 396.000 83.630 400.000 ;
    END
  END dout0_to_sram[13]
  PIN dout0_to_sram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END dout0_to_sram[14]
  PIN dout0_to_sram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 396.000 96.050 400.000 ;
    END
  END dout0_to_sram[15]
  PIN dout0_to_sram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END dout0_to_sram[16]
  PIN dout0_to_sram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.240 400.000 112.840 ;
    END
  END dout0_to_sram[17]
  PIN dout0_to_sram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END dout0_to_sram[18]
  PIN dout0_to_sram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END dout0_to_sram[19]
  PIN dout0_to_sram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END dout0_to_sram[1]
  PIN dout0_to_sram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 396.000 132.390 400.000 ;
    END
  END dout0_to_sram[20]
  PIN dout0_to_sram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 396.000 135.610 400.000 ;
    END
  END dout0_to_sram[21]
  PIN dout0_to_sram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 396.000 144.350 400.000 ;
    END
  END dout0_to_sram[22]
  PIN dout0_to_sram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END dout0_to_sram[23]
  PIN dout0_to_sram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 154.400 400.000 155.000 ;
    END
  END dout0_to_sram[24]
  PIN dout0_to_sram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 396.000 158.150 400.000 ;
    END
  END dout0_to_sram[25]
  PIN dout0_to_sram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 165.280 400.000 165.880 ;
    END
  END dout0_to_sram[26]
  PIN dout0_to_sram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END dout0_to_sram[27]
  PIN dout0_to_sram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END dout0_to_sram[28]
  PIN dout0_to_sram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END dout0_to_sram[29]
  PIN dout0_to_sram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END dout0_to_sram[2]
  PIN dout0_to_sram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END dout0_to_sram[30]
  PIN dout0_to_sram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END dout0_to_sram[31]
  PIN dout0_to_sram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END dout0_to_sram[3]
  PIN dout0_to_sram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 32.680 400.000 33.280 ;
    END
  END dout0_to_sram[4]
  PIN dout0_to_sram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END dout0_to_sram[5]
  PIN dout0_to_sram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END dout0_to_sram[6]
  PIN dout0_to_sram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 396.000 42.230 400.000 ;
    END
  END dout0_to_sram[7]
  PIN dout0_to_sram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 65.320 400.000 65.920 ;
    END
  END dout0_to_sram[8]
  PIN dout0_to_sram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 70.080 400.000 70.680 ;
    END
  END dout0_to_sram[9]
  PIN is_loading_memory_into_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END is_loading_memory_into_core
  PIN is_ready_dataout_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END is_ready_dataout_core0
  PIN is_ready_print_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END is_ready_print_core0
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 396.000 340.310 400.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 343.440 400.000 344.040 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 74.840 400.000 75.440 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 396.000 364.230 400.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 396.000 366.070 400.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 396.000 369.750 400.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 369.280 400.000 369.880 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 372.680 400.000 373.280 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 396.000 381.710 400.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 396.000 390.450 400.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 379.480 400.000 380.080 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 396.000 395.510 400.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 384.240 400.000 384.840 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 389.000 400.000 389.600 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 395.120 400.000 395.720 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 87.760 400.000 88.360 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 99.320 400.000 99.920 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 113.600 400.000 114.200 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 118.360 400.000 118.960 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.920 400.000 130.520 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 131.280 400.000 131.880 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 396.000 137.450 400.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 146.240 400.000 146.840 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 155.760 400.000 156.360 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 396.000 170.570 400.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 396.000 178.850 400.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 18.400 400.000 19.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 181.600 400.000 182.200 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 196.560 400.000 197.160 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 396.000 196.330 400.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 201.320 400.000 201.920 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 202.680 400.000 203.280 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 396.000 208.290 400.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 212.200 400.000 212.800 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.960 400.000 217.560 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 396.000 218.870 400.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 225.120 400.000 225.720 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 34.040 400.000 34.640 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 396.000 225.770 400.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 240.080 400.000 240.680 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 396.000 236.350 400.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 396.000 243.250 400.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 396.000 248.310 400.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 261.160 400.000 261.760 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 396.000 262.110 400.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 396.000 267.630 400.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.840 400.000 279.440 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 396.000 275.910 400.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 288.360 400.000 288.960 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 396.000 288.330 400.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 293.120 400.000 293.720 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 296.520 400.000 297.120 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 396.000 307.190 400.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 298.560 400.000 299.160 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.040 400.000 306.640 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 396.000 315.930 400.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 396.000 317.770 400.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 312.840 400.000 313.440 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 396.000 320.990 400.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 396.000 326.510 400.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 396.000 327.890 400.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 324.400 400.000 325.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 327.120 400.000 327.720 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 396.000 0.830 400.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 335.280 400.000 335.880 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 340.040 400.000 340.640 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 396.000 341.690 400.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 396.000 349.050 400.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 352.960 400.000 353.560 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 396.000 355.950 400.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 396.000 357.330 400.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 396.000 361.010 400.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 363.160 400.000 363.760 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 396.000 367.910 400.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 371.320 400.000 371.920 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 396.000 376.650 400.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 396.000 383.550 400.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 396.000 397.350 400.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 396.000 399.190 400.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 390.360 400.000 390.960 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 89.120 400.000 89.720 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 396.000 97.430 400.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 396.000 106.170 400.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 396.000 113.070 400.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 396.000 10.950 400.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 160.520 400.000 161.120 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 396.000 171.950 400.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 396.000 180.690 400.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 396.000 185.750 400.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 396.000 21.530 400.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 185.000 400.000 185.600 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 191.120 400.000 191.720 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 199.280 400.000 199.880 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 396.000 203.230 400.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.040 400.000 204.640 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 209.480 400.000 210.080 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 396.000 211.970 400.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 396.000 213.810 400.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 215.600 400.000 216.200 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 222.400 400.000 223.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 396.000 223.930 400.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 230.560 400.000 231.160 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 36.080 400.000 36.680 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.040 400.000 238.640 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 396.000 237.730 400.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.240 400.000 248.840 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 253.000 400.000 253.600 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 47.640 400.000 48.240 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 257.760 400.000 258.360 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 396.000 255.210 400.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 264.560 400.000 265.160 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 267.280 400.000 267.880 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 272.040 400.000 272.640 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 282.240 400.000 282.840 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 396.000 272.690 400.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 396.000 279.590 400.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 290.400 400.000 291.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 396.000 289.710 400.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 396.000 295.230 400.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 396.000 303.970 400.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 301.280 400.000 301.880 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 4.000 325.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 309.440 400.000 310.040 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 396.000 319.150 400.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 396.000 329.730 400.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 396.000 334.790 400.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 329.160 400.000 329.760 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 396.000 59.710 400.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 396.000 2.210 400.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 396.000 336.630 400.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 396.000 343.530 400.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 396.000 345.370 400.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 346.840 400.000 347.440 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 348.200 400.000 348.800 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 351.600 400.000 352.200 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 396.000 354.110 400.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 356.360 400.000 356.960 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 359.760 400.000 360.360 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 396.000 371.130 400.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 367.920 400.000 368.520 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 396.000 378.490 400.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 396.000 71.670 400.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 376.080 400.000 376.680 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 380.840 400.000 381.440 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 385.600 400.000 386.200 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 393.760 400.000 394.360 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 397.160 400.000 397.760 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 396.000 123.650 400.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 11.600 400.000 12.200 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 138.080 400.000 138.680 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 396.000 146.190 400.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 147.600 400.000 148.200 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 396.000 153.090 400.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 396.000 173.790 400.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 396.000 187.590 400.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 396.000 22.910 400.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 186.360 400.000 186.960 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.160 400.000 193.760 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.920 400.000 198.520 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 396.000 198.170 400.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 396.000 205.070 400.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 206.080 400.000 206.680 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 396.000 206.910 400.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 396.000 26.590 400.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 396.000 215.650 400.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 219.000 400.000 219.600 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 396.000 220.710 400.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.160 400.000 227.760 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 231.920 400.000 232.520 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 37.440 400.000 38.040 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 396.000 227.610 400.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 396.000 230.830 400.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 241.440 400.000 242.040 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 396.000 239.570 400.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 244.840 400.000 245.440 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 249.600 400.000 250.200 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 396.000 246.470 400.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 259.120 400.000 259.720 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 396.000 251.990 400.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 396.000 257.050 400.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 262.520 400.000 263.120 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 396.000 263.950 400.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 55.120 400.000 55.720 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 275.440 400.000 276.040 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 280.200 400.000 280.800 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 283.600 400.000 284.200 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 284.960 400.000 285.560 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 396.000 277.750 400.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 396.000 281.430 400.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 396.000 284.650 400.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 396.000 44.070 400.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 291.760 400.000 292.360 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 396.000 297.070 400.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 295.160 400.000 295.760 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 396.000 305.350 400.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 396.000 309.030 400.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 304.680 400.000 305.280 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 396.000 314.090 400.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 396.000 52.350 400.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 396.000 322.830 400.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 317.600 400.000 318.200 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 396.000 331.570 400.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END la_oenb[9]
  PIN rd_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END rd_data_out[0]
  PIN rd_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 332.560 400.000 333.160 ;
    END
  END rd_data_out[100]
  PIN rd_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 337.320 400.000 337.920 ;
    END
  END rd_data_out[101]
  PIN rd_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 396.000 338.470 400.000 ;
    END
  END rd_data_out[102]
  PIN rd_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END rd_data_out[103]
  PIN rd_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 345.480 400.000 346.080 ;
    END
  END rd_data_out[104]
  PIN rd_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END rd_data_out[105]
  PIN rd_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 396.000 350.430 400.000 ;
    END
  END rd_data_out[106]
  PIN rd_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END rd_data_out[107]
  PIN rd_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END rd_data_out[108]
  PIN rd_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 355.000 400.000 355.600 ;
    END
  END rd_data_out[109]
  PIN rd_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 396.000 64.770 400.000 ;
    END
  END rd_data_out[10]
  PIN rd_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END rd_data_out[110]
  PIN rd_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 396.000 359.170 400.000 ;
    END
  END rd_data_out[111]
  PIN rd_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 361.120 400.000 361.720 ;
    END
  END rd_data_out[112]
  PIN rd_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 364.520 400.000 365.120 ;
    END
  END rd_data_out[113]
  PIN rd_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END rd_data_out[114]
  PIN rd_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 366.560 400.000 367.160 ;
    END
  END rd_data_out[115]
  PIN rd_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 396.000 374.810 400.000 ;
    END
  END rd_data_out[116]
  PIN rd_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END rd_data_out[117]
  PIN rd_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 396.000 379.870 400.000 ;
    END
  END rd_data_out[118]
  PIN rd_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 396.000 385.390 400.000 ;
    END
  END rd_data_out[119]
  PIN rd_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END rd_data_out[11]
  PIN rd_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 396.000 386.770 400.000 ;
    END
  END rd_data_out[120]
  PIN rd_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 377.440 400.000 378.040 ;
    END
  END rd_data_out[121]
  PIN rd_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 396.000 392.290 400.000 ;
    END
  END rd_data_out[122]
  PIN rd_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 382.200 400.000 382.800 ;
    END
  END rd_data_out[123]
  PIN rd_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 386.960 400.000 387.560 ;
    END
  END rd_data_out[124]
  PIN rd_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 392.400 400.000 393.000 ;
    END
  END rd_data_out[125]
  PIN rd_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END rd_data_out[126]
  PIN rd_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 398.520 400.000 399.120 ;
    END
  END rd_data_out[127]
  PIN rd_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END rd_data_out[12]
  PIN rd_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END rd_data_out[13]
  PIN rd_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END rd_data_out[14]
  PIN rd_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END rd_data_out[15]
  PIN rd_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END rd_data_out[16]
  PIN rd_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 115.640 400.000 116.240 ;
    END
  END rd_data_out[17]
  PIN rd_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 120.400 400.000 121.000 ;
    END
  END rd_data_out[18]
  PIN rd_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 396.000 126.870 400.000 ;
    END
  END rd_data_out[19]
  PIN rd_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 13.640 400.000 14.240 ;
    END
  END rd_data_out[1]
  PIN rd_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END rd_data_out[20]
  PIN rd_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END rd_data_out[21]
  PIN rd_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 396.000 148.030 400.000 ;
    END
  END rd_data_out[22]
  PIN rd_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 149.640 400.000 150.240 ;
    END
  END rd_data_out[23]
  PIN rd_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END rd_data_out[24]
  PIN rd_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 162.560 400.000 163.160 ;
    END
  END rd_data_out[25]
  PIN rd_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 167.320 400.000 167.920 ;
    END
  END rd_data_out[26]
  PIN rd_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.040 400.000 170.640 ;
    END
  END rd_data_out[27]
  PIN rd_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END rd_data_out[28]
  PIN rd_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END rd_data_out[29]
  PIN rd_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 396.000 24.750 400.000 ;
    END
  END rd_data_out[2]
  PIN rd_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END rd_data_out[30]
  PIN rd_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 188.400 400.000 189.000 ;
    END
  END rd_data_out[31]
  PIN rd_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 194.520 400.000 195.120 ;
    END
  END rd_data_out[32]
  PIN rd_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END rd_data_out[33]
  PIN rd_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 396.000 193.110 400.000 ;
    END
  END rd_data_out[34]
  PIN rd_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 396.000 200.010 400.000 ;
    END
  END rd_data_out[35]
  PIN rd_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END rd_data_out[36]
  PIN rd_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END rd_data_out[37]
  PIN rd_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END rd_data_out[38]
  PIN rd_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END rd_data_out[39]
  PIN rd_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 396.000 28.430 400.000 ;
    END
  END rd_data_out[3]
  PIN rd_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.840 400.000 211.440 ;
    END
  END rd_data_out[40]
  PIN rd_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END rd_data_out[41]
  PIN rd_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END rd_data_out[42]
  PIN rd_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END rd_data_out[43]
  PIN rd_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END rd_data_out[44]
  PIN rd_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 220.360 400.000 220.960 ;
    END
  END rd_data_out[45]
  PIN rd_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 396.000 222.550 400.000 ;
    END
  END rd_data_out[46]
  PIN rd_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 228.520 400.000 229.120 ;
    END
  END rd_data_out[47]
  PIN rd_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END rd_data_out[48]
  PIN rd_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 233.280 400.000 233.880 ;
    END
  END rd_data_out[49]
  PIN rd_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 396.000 31.650 400.000 ;
    END
  END rd_data_out[4]
  PIN rd_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END rd_data_out[50]
  PIN rd_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END rd_data_out[51]
  PIN rd_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 396.000 229.450 400.000 ;
    END
  END rd_data_out[52]
  PIN rd_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END rd_data_out[53]
  PIN rd_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 396.000 232.670 400.000 ;
    END
  END rd_data_out[54]
  PIN rd_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 243.480 400.000 244.080 ;
    END
  END rd_data_out[55]
  PIN rd_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 396.000 241.410 400.000 ;
    END
  END rd_data_out[56]
  PIN rd_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END rd_data_out[57]
  PIN rd_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 396.000 245.090 400.000 ;
    END
  END rd_data_out[58]
  PIN rd_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 254.360 400.000 254.960 ;
    END
  END rd_data_out[59]
  PIN rd_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END rd_data_out[5]
  PIN rd_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END rd_data_out[60]
  PIN rd_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 256.400 400.000 257.000 ;
    END
  END rd_data_out[61]
  PIN rd_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END rd_data_out[62]
  PIN rd_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 396.000 253.370 400.000 ;
    END
  END rd_data_out[63]
  PIN rd_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END rd_data_out[64]
  PIN rd_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END rd_data_out[65]
  PIN rd_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END rd_data_out[66]
  PIN rd_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 396.000 260.270 400.000 ;
    END
  END rd_data_out[67]
  PIN rd_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END rd_data_out[68]
  PIN rd_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 396.000 265.790 400.000 ;
    END
  END rd_data_out[69]
  PIN rd_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END rd_data_out[6]
  PIN rd_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 269.320 400.000 269.920 ;
    END
  END rd_data_out[70]
  PIN rd_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 274.080 400.000 274.680 ;
    END
  END rd_data_out[71]
  PIN rd_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 277.480 400.000 278.080 ;
    END
  END rd_data_out[72]
  PIN rd_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END rd_data_out[73]
  PIN rd_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 396.000 269.010 400.000 ;
    END
  END rd_data_out[74]
  PIN rd_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 396.000 274.530 400.000 ;
    END
  END rd_data_out[75]
  PIN rd_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END rd_data_out[76]
  PIN rd_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 396.000 282.810 400.000 ;
    END
  END rd_data_out[77]
  PIN rd_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END rd_data_out[78]
  PIN rd_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END rd_data_out[79]
  PIN rd_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 396.000 45.450 400.000 ;
    END
  END rd_data_out[7]
  PIN rd_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 396.000 293.390 400.000 ;
    END
  END rd_data_out[80]
  PIN rd_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 396.000 298.450 400.000 ;
    END
  END rd_data_out[81]
  PIN rd_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END rd_data_out[82]
  PIN rd_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END rd_data_out[83]
  PIN rd_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END rd_data_out[84]
  PIN rd_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 299.920 400.000 300.520 ;
    END
  END rd_data_out[85]
  PIN rd_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 303.320 400.000 303.920 ;
    END
  END rd_data_out[86]
  PIN rd_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 396.000 312.250 400.000 ;
    END
  END rd_data_out[87]
  PIN rd_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END rd_data_out[88]
  PIN rd_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END rd_data_out[89]
  PIN rd_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 396.000 54.190 400.000 ;
    END
  END rd_data_out[8]
  PIN rd_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 311.480 400.000 312.080 ;
    END
  END rd_data_out[90]
  PIN rd_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 314.200 400.000 314.800 ;
    END
  END rd_data_out[91]
  PIN rd_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END rd_data_out[92]
  PIN rd_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 318.960 400.000 319.560 ;
    END
  END rd_data_out[93]
  PIN rd_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.000 400.000 321.600 ;
    END
  END rd_data_out[94]
  PIN rd_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END rd_data_out[95]
  PIN rd_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END rd_data_out[96]
  PIN rd_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 396.000 333.410 400.000 ;
    END
  END rd_data_out[97]
  PIN rd_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 325.760 400.000 326.360 ;
    END
  END rd_data_out[98]
  PIN rd_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END rd_data_out[99]
  PIN rd_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END rd_data_out[9]
  PIN read_enable_to_Elpis
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END read_enable_to_Elpis
  PIN read_interactive_req_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END read_interactive_req_core0
  PIN read_value_to_Elpis[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 396.000 4.050 400.000 ;
    END
  END read_value_to_Elpis[0]
  PIN read_value_to_Elpis[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 396.000 66.610 400.000 ;
    END
  END read_value_to_Elpis[10]
  PIN read_value_to_Elpis[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 81.640 400.000 82.240 ;
    END
  END read_value_to_Elpis[11]
  PIN read_value_to_Elpis[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 396.000 76.730 400.000 ;
    END
  END read_value_to_Elpis[12]
  PIN read_value_to_Elpis[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 91.160 400.000 91.760 ;
    END
  END read_value_to_Elpis[13]
  PIN read_value_to_Elpis[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 396.000 90.530 400.000 ;
    END
  END read_value_to_Elpis[14]
  PIN read_value_to_Elpis[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 100.680 400.000 101.280 ;
    END
  END read_value_to_Elpis[15]
  PIN read_value_to_Elpis[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 105.440 400.000 106.040 ;
    END
  END read_value_to_Elpis[16]
  PIN read_value_to_Elpis[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 396.000 114.910 400.000 ;
    END
  END read_value_to_Elpis[17]
  PIN read_value_to_Elpis[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 121.760 400.000 122.360 ;
    END
  END read_value_to_Elpis[18]
  PIN read_value_to_Elpis[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END read_value_to_Elpis[19]
  PIN read_value_to_Elpis[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 15.000 400.000 15.600 ;
    END
  END read_value_to_Elpis[1]
  PIN read_value_to_Elpis[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END read_value_to_Elpis[20]
  PIN read_value_to_Elpis[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 396.000 139.290 400.000 ;
    END
  END read_value_to_Elpis[21]
  PIN read_value_to_Elpis[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 396.000 149.410 400.000 ;
    END
  END read_value_to_Elpis[22]
  PIN read_value_to_Elpis[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 151.000 400.000 151.600 ;
    END
  END read_value_to_Elpis[23]
  PIN read_value_to_Elpis[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END read_value_to_Elpis[24]
  PIN read_value_to_Elpis[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 396.000 159.990 400.000 ;
    END
  END read_value_to_Elpis[25]
  PIN read_value_to_Elpis[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 396.000 166.890 400.000 ;
    END
  END read_value_to_Elpis[26]
  PIN read_value_to_Elpis[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 396.000 175.630 400.000 ;
    END
  END read_value_to_Elpis[27]
  PIN read_value_to_Elpis[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 396.000 182.530 400.000 ;
    END
  END read_value_to_Elpis[28]
  PIN read_value_to_Elpis[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END read_value_to_Elpis[29]
  PIN read_value_to_Elpis[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 19.760 400.000 20.360 ;
    END
  END read_value_to_Elpis[2]
  PIN read_value_to_Elpis[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END read_value_to_Elpis[30]
  PIN read_value_to_Elpis[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END read_value_to_Elpis[31]
  PIN read_value_to_Elpis[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END read_value_to_Elpis[3]
  PIN read_value_to_Elpis[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END read_value_to_Elpis[4]
  PIN read_value_to_Elpis[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 49.000 400.000 49.600 ;
    END
  END read_value_to_Elpis[5]
  PIN read_value_to_Elpis[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 396.000 38.550 400.000 ;
    END
  END read_value_to_Elpis[6]
  PIN read_value_to_Elpis[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 60.560 400.000 61.160 ;
    END
  END read_value_to_Elpis[7]
  PIN read_value_to_Elpis[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END read_value_to_Elpis[8]
  PIN read_value_to_Elpis[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 71.440 400.000 72.040 ;
    END
  END read_value_to_Elpis[9]
  PIN ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END ready
  PIN req_out_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END req_out_core0
  PIN requested
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END requested
  PIN reset_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END reset_core
  PIN reset_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END reset_mem_req
  PIN rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END rst
  PIN spare_wen0_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 3.440 400.000 4.040 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_rst_i
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 396.000 5.890 400.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 396.000 73.510 400.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 396.000 85.470 400.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.920 400.000 96.520 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 396.000 99.270 400.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 396.000 108.010 400.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 396.000 128.710 400.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 16.360 400.000 16.960 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 133.320 400.000 133.920 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 139.440 400.000 140.040 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 141.480 400.000 142.080 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 157.120 400.000 157.720 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 172.080 400.000 172.680 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 396.000 184.370 400.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 178.200 400.000 178.800 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 396.000 33.490 400.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 396.000 37.170 400.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 61.920 400.000 62.520 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 396.000 56.030 400.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 396.000 61.090 400.000 ;
    END
  END wbs_dat_o[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END we
  PIN we_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 0.720 400.000 1.320 ;
    END
  END we_to_sram
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 396.000 7.730 400.000 ;
    END
  END wr_data[0]
  PIN wr_data[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.920 400.000 334.520 ;
    END
  END wr_data[100]
  PIN wr_data[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 338.680 400.000 339.280 ;
    END
  END wr_data[101]
  PIN wr_data[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END wr_data[102]
  PIN wr_data[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 342.080 400.000 342.680 ;
    END
  END wr_data[103]
  PIN wr_data[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 396.000 347.210 400.000 ;
    END
  END wr_data[104]
  PIN wr_data[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END wr_data[105]
  PIN wr_data[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END wr_data[106]
  PIN wr_data[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 350.240 400.000 350.840 ;
    END
  END wr_data[107]
  PIN wr_data[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 396.000 352.270 400.000 ;
    END
  END wr_data[108]
  PIN wr_data[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END wr_data[109]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 76.200 400.000 76.800 ;
    END
  END wr_data[10]
  PIN wr_data[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END wr_data[110]
  PIN wr_data[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 358.400 400.000 359.000 ;
    END
  END wr_data[111]
  PIN wr_data[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 396.000 362.850 400.000 ;
    END
  END wr_data[112]
  PIN wr_data[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END wr_data[113]
  PIN wr_data[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END wr_data[114]
  PIN wr_data[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 396.000 372.970 400.000 ;
    END
  END wr_data[115]
  PIN wr_data[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END wr_data[116]
  PIN wr_data[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END wr_data[117]
  PIN wr_data[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END wr_data[118]
  PIN wr_data[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 374.040 400.000 374.640 ;
    END
  END wr_data[119]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END wr_data[11]
  PIN wr_data[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 396.000 388.610 400.000 ;
    END
  END wr_data[120]
  PIN wr_data[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END wr_data[121]
  PIN wr_data[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 396.000 393.670 400.000 ;
    END
  END wr_data[122]
  PIN wr_data[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END wr_data[123]
  PIN wr_data[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END wr_data[124]
  PIN wr_data[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END wr_data[125]
  PIN wr_data[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END wr_data[126]
  PIN wr_data[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END wr_data[127]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 86.400 400.000 87.000 ;
    END
  END wr_data[12]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END wr_data[13]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wr_data[14]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wr_data[15]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 396.000 109.850 400.000 ;
    END
  END wr_data[16]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 396.000 116.750 400.000 ;
    END
  END wr_data[17]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 396.000 125.490 400.000 ;
    END
  END wr_data[18]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 396.000 130.550 400.000 ;
    END
  END wr_data[19]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 396.000 12.790 400.000 ;
    END
  END wr_data[1]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 396.000 134.230 400.000 ;
    END
  END wr_data[20]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wr_data[21]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 396.000 151.250 400.000 ;
    END
  END wr_data[22]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 152.360 400.000 152.960 ;
    END
  END wr_data[23]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END wr_data[24]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 396.000 161.830 400.000 ;
    END
  END wr_data[25]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 396.000 168.730 400.000 ;
    END
  END wr_data[26]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 173.440 400.000 174.040 ;
    END
  END wr_data[27]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END wr_data[28]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 396.000 189.430 400.000 ;
    END
  END wr_data[29]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END wr_data[2]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 396.000 191.270 400.000 ;
    END
  END wr_data[30]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 189.760 400.000 190.360 ;
    END
  END wr_data[31]
  PIN wr_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END wr_data[32]
  PIN wr_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END wr_data[33]
  PIN wr_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 396.000 194.490 400.000 ;
    END
  END wr_data[34]
  PIN wr_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 396.000 201.390 400.000 ;
    END
  END wr_data[35]
  PIN wr_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END wr_data[36]
  PIN wr_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END wr_data[37]
  PIN wr_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 207.440 400.000 208.040 ;
    END
  END wr_data[38]
  PIN wr_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wr_data[39]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 396.000 30.270 400.000 ;
    END
  END wr_data[3]
  PIN wr_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 396.000 210.130 400.000 ;
    END
  END wr_data[40]
  PIN wr_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END wr_data[41]
  PIN wr_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.240 400.000 214.840 ;
    END
  END wr_data[42]
  PIN wr_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 396.000 217.030 400.000 ;
    END
  END wr_data[43]
  PIN wr_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END wr_data[44]
  PIN wr_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wr_data[45]
  PIN wr_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 223.760 400.000 224.360 ;
    END
  END wr_data[46]
  PIN wr_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wr_data[47]
  PIN wr_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END wr_data[48]
  PIN wr_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END wr_data[49]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 396.000 35.330 400.000 ;
    END
  END wr_data[4]
  PIN wr_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 235.320 400.000 235.920 ;
    END
  END wr_data[50]
  PIN wr_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 236.680 400.000 237.280 ;
    END
  END wr_data[51]
  PIN wr_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END wr_data[52]
  PIN wr_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END wr_data[53]
  PIN wr_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 396.000 234.510 400.000 ;
    END
  END wr_data[54]
  PIN wr_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END wr_data[55]
  PIN wr_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END wr_data[56]
  PIN wr_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 246.200 400.000 246.800 ;
    END
  END wr_data[57]
  PIN wr_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 250.960 400.000 251.560 ;
    END
  END wr_data[58]
  PIN wr_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END wr_data[59]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END wr_data[5]
  PIN wr_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wr_data[60]
  PIN wr_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 396.000 250.150 400.000 ;
    END
  END wr_data[61]
  PIN wr_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END wr_data[62]
  PIN wr_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wr_data[63]
  PIN wr_data[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wr_data[64]
  PIN wr_data[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wr_data[65]
  PIN wr_data[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 396.000 258.890 400.000 ;
    END
  END wr_data[66]
  PIN wr_data[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END wr_data[67]
  PIN wr_data[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END wr_data[68]
  PIN wr_data[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.920 400.000 266.520 ;
    END
  END wr_data[69]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 57.160 400.000 57.760 ;
    END
  END wr_data[6]
  PIN wr_data[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 270.680 400.000 271.280 ;
    END
  END wr_data[70]
  PIN wr_data[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END wr_data[71]
  PIN wr_data[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END wr_data[72]
  PIN wr_data[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END wr_data[73]
  PIN wr_data[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 396.000 270.850 400.000 ;
    END
  END wr_data[74]
  PIN wr_data[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 287.000 400.000 287.600 ;
    END
  END wr_data[75]
  PIN wr_data[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END wr_data[76]
  PIN wr_data[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wr_data[77]
  PIN wr_data[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 396.000 286.490 400.000 ;
    END
  END wr_data[78]
  PIN wr_data[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 396.000 291.550 400.000 ;
    END
  END wr_data[79]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END wr_data[7]
  PIN wr_data[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END wr_data[80]
  PIN wr_data[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 396.000 300.290 400.000 ;
    END
  END wr_data[81]
  PIN wr_data[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 396.000 302.130 400.000 ;
    END
  END wr_data[82]
  PIN wr_data[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END wr_data[83]
  PIN wr_data[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END wr_data[84]
  PIN wr_data[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END wr_data[85]
  PIN wr_data[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 396.000 310.870 400.000 ;
    END
  END wr_data[86]
  PIN wr_data[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END wr_data[87]
  PIN wr_data[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 308.080 400.000 308.680 ;
    END
  END wr_data[88]
  PIN wr_data[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END wr_data[89]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END wr_data[8]
  PIN wr_data[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END wr_data[90]
  PIN wr_data[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 316.240 400.000 316.840 ;
    END
  END wr_data[91]
  PIN wr_data[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END wr_data[92]
  PIN wr_data[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END wr_data[93]
  PIN wr_data[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 396.000 324.670 400.000 ;
    END
  END wr_data[94]
  PIN wr_data[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END wr_data[95]
  PIN wr_data[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 322.360 400.000 322.960 ;
    END
  END wr_data[96]
  PIN wr_data[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END wr_data[97]
  PIN wr_data[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END wr_data[98]
  PIN wr_data[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 330.520 400.000 331.120 ;
    END
  END wr_data[99]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wr_data[9]
  OBS
      LAYER li1 ;
        RECT 5.520 7.225 396.835 391.935 ;
      LAYER met1 ;
        RECT 0.530 4.460 399.210 393.000 ;
      LAYER met2 ;
        RECT 1.110 395.720 1.650 399.005 ;
        RECT 2.490 395.720 3.490 399.005 ;
        RECT 4.330 395.720 5.330 399.005 ;
        RECT 6.170 395.720 7.170 399.005 ;
        RECT 8.010 395.720 8.550 399.005 ;
        RECT 9.390 395.720 10.390 399.005 ;
        RECT 11.230 395.720 12.230 399.005 ;
        RECT 13.070 395.720 14.070 399.005 ;
        RECT 14.910 395.720 15.450 399.005 ;
        RECT 16.290 395.720 17.290 399.005 ;
        RECT 18.130 395.720 19.130 399.005 ;
        RECT 19.970 395.720 20.970 399.005 ;
        RECT 21.810 395.720 22.350 399.005 ;
        RECT 23.190 395.720 24.190 399.005 ;
        RECT 25.030 395.720 26.030 399.005 ;
        RECT 26.870 395.720 27.870 399.005 ;
        RECT 28.710 395.720 29.710 399.005 ;
        RECT 30.550 395.720 31.090 399.005 ;
        RECT 31.930 395.720 32.930 399.005 ;
        RECT 33.770 395.720 34.770 399.005 ;
        RECT 35.610 395.720 36.610 399.005 ;
        RECT 37.450 395.720 37.990 399.005 ;
        RECT 38.830 395.720 39.830 399.005 ;
        RECT 40.670 395.720 41.670 399.005 ;
        RECT 42.510 395.720 43.510 399.005 ;
        RECT 44.350 395.720 44.890 399.005 ;
        RECT 45.730 395.720 46.730 399.005 ;
        RECT 47.570 395.720 48.570 399.005 ;
        RECT 49.410 395.720 50.410 399.005 ;
        RECT 51.250 395.720 51.790 399.005 ;
        RECT 52.630 395.720 53.630 399.005 ;
        RECT 54.470 395.720 55.470 399.005 ;
        RECT 56.310 395.720 57.310 399.005 ;
        RECT 58.150 395.720 59.150 399.005 ;
        RECT 59.990 395.720 60.530 399.005 ;
        RECT 61.370 395.720 62.370 399.005 ;
        RECT 63.210 395.720 64.210 399.005 ;
        RECT 65.050 395.720 66.050 399.005 ;
        RECT 66.890 395.720 67.430 399.005 ;
        RECT 68.270 395.720 69.270 399.005 ;
        RECT 70.110 395.720 71.110 399.005 ;
        RECT 71.950 395.720 72.950 399.005 ;
        RECT 73.790 395.720 74.330 399.005 ;
        RECT 75.170 395.720 76.170 399.005 ;
        RECT 77.010 395.720 78.010 399.005 ;
        RECT 78.850 395.720 79.850 399.005 ;
        RECT 80.690 395.720 81.690 399.005 ;
        RECT 82.530 395.720 83.070 399.005 ;
        RECT 83.910 395.720 84.910 399.005 ;
        RECT 85.750 395.720 86.750 399.005 ;
        RECT 87.590 395.720 88.590 399.005 ;
        RECT 89.430 395.720 89.970 399.005 ;
        RECT 90.810 395.720 91.810 399.005 ;
        RECT 92.650 395.720 93.650 399.005 ;
        RECT 94.490 395.720 95.490 399.005 ;
        RECT 96.330 395.720 96.870 399.005 ;
        RECT 97.710 395.720 98.710 399.005 ;
        RECT 99.550 395.720 100.550 399.005 ;
        RECT 101.390 395.720 102.390 399.005 ;
        RECT 103.230 395.720 103.770 399.005 ;
        RECT 104.610 395.720 105.610 399.005 ;
        RECT 106.450 395.720 107.450 399.005 ;
        RECT 108.290 395.720 109.290 399.005 ;
        RECT 110.130 395.720 111.130 399.005 ;
        RECT 111.970 395.720 112.510 399.005 ;
        RECT 113.350 395.720 114.350 399.005 ;
        RECT 115.190 395.720 116.190 399.005 ;
        RECT 117.030 395.720 118.030 399.005 ;
        RECT 118.870 395.720 119.410 399.005 ;
        RECT 120.250 395.720 121.250 399.005 ;
        RECT 122.090 395.720 123.090 399.005 ;
        RECT 123.930 395.720 124.930 399.005 ;
        RECT 125.770 395.720 126.310 399.005 ;
        RECT 127.150 395.720 128.150 399.005 ;
        RECT 128.990 395.720 129.990 399.005 ;
        RECT 130.830 395.720 131.830 399.005 ;
        RECT 132.670 395.720 133.670 399.005 ;
        RECT 134.510 395.720 135.050 399.005 ;
        RECT 135.890 395.720 136.890 399.005 ;
        RECT 137.730 395.720 138.730 399.005 ;
        RECT 139.570 395.720 140.570 399.005 ;
        RECT 141.410 395.720 141.950 399.005 ;
        RECT 142.790 395.720 143.790 399.005 ;
        RECT 144.630 395.720 145.630 399.005 ;
        RECT 146.470 395.720 147.470 399.005 ;
        RECT 148.310 395.720 148.850 399.005 ;
        RECT 149.690 395.720 150.690 399.005 ;
        RECT 151.530 395.720 152.530 399.005 ;
        RECT 153.370 395.720 154.370 399.005 ;
        RECT 155.210 395.720 155.750 399.005 ;
        RECT 156.590 395.720 157.590 399.005 ;
        RECT 158.430 395.720 159.430 399.005 ;
        RECT 160.270 395.720 161.270 399.005 ;
        RECT 162.110 395.720 163.110 399.005 ;
        RECT 163.950 395.720 164.490 399.005 ;
        RECT 165.330 395.720 166.330 399.005 ;
        RECT 167.170 395.720 168.170 399.005 ;
        RECT 169.010 395.720 170.010 399.005 ;
        RECT 170.850 395.720 171.390 399.005 ;
        RECT 172.230 395.720 173.230 399.005 ;
        RECT 174.070 395.720 175.070 399.005 ;
        RECT 175.910 395.720 176.910 399.005 ;
        RECT 177.750 395.720 178.290 399.005 ;
        RECT 179.130 395.720 180.130 399.005 ;
        RECT 180.970 395.720 181.970 399.005 ;
        RECT 182.810 395.720 183.810 399.005 ;
        RECT 184.650 395.720 185.190 399.005 ;
        RECT 186.030 395.720 187.030 399.005 ;
        RECT 187.870 395.720 188.870 399.005 ;
        RECT 189.710 395.720 190.710 399.005 ;
        RECT 191.550 395.720 192.550 399.005 ;
        RECT 193.390 395.720 193.930 399.005 ;
        RECT 194.770 395.720 195.770 399.005 ;
        RECT 196.610 395.720 197.610 399.005 ;
        RECT 198.450 395.720 199.450 399.005 ;
        RECT 200.290 395.720 200.830 399.005 ;
        RECT 201.670 395.720 202.670 399.005 ;
        RECT 203.510 395.720 204.510 399.005 ;
        RECT 205.350 395.720 206.350 399.005 ;
        RECT 207.190 395.720 207.730 399.005 ;
        RECT 208.570 395.720 209.570 399.005 ;
        RECT 210.410 395.720 211.410 399.005 ;
        RECT 212.250 395.720 213.250 399.005 ;
        RECT 214.090 395.720 215.090 399.005 ;
        RECT 215.930 395.720 216.470 399.005 ;
        RECT 217.310 395.720 218.310 399.005 ;
        RECT 219.150 395.720 220.150 399.005 ;
        RECT 220.990 395.720 221.990 399.005 ;
        RECT 222.830 395.720 223.370 399.005 ;
        RECT 224.210 395.720 225.210 399.005 ;
        RECT 226.050 395.720 227.050 399.005 ;
        RECT 227.890 395.720 228.890 399.005 ;
        RECT 229.730 395.720 230.270 399.005 ;
        RECT 231.110 395.720 232.110 399.005 ;
        RECT 232.950 395.720 233.950 399.005 ;
        RECT 234.790 395.720 235.790 399.005 ;
        RECT 236.630 395.720 237.170 399.005 ;
        RECT 238.010 395.720 239.010 399.005 ;
        RECT 239.850 395.720 240.850 399.005 ;
        RECT 241.690 395.720 242.690 399.005 ;
        RECT 243.530 395.720 244.530 399.005 ;
        RECT 245.370 395.720 245.910 399.005 ;
        RECT 246.750 395.720 247.750 399.005 ;
        RECT 248.590 395.720 249.590 399.005 ;
        RECT 250.430 395.720 251.430 399.005 ;
        RECT 252.270 395.720 252.810 399.005 ;
        RECT 253.650 395.720 254.650 399.005 ;
        RECT 255.490 395.720 256.490 399.005 ;
        RECT 257.330 395.720 258.330 399.005 ;
        RECT 259.170 395.720 259.710 399.005 ;
        RECT 260.550 395.720 261.550 399.005 ;
        RECT 262.390 395.720 263.390 399.005 ;
        RECT 264.230 395.720 265.230 399.005 ;
        RECT 266.070 395.720 267.070 399.005 ;
        RECT 267.910 395.720 268.450 399.005 ;
        RECT 269.290 395.720 270.290 399.005 ;
        RECT 271.130 395.720 272.130 399.005 ;
        RECT 272.970 395.720 273.970 399.005 ;
        RECT 274.810 395.720 275.350 399.005 ;
        RECT 276.190 395.720 277.190 399.005 ;
        RECT 278.030 395.720 279.030 399.005 ;
        RECT 279.870 395.720 280.870 399.005 ;
        RECT 281.710 395.720 282.250 399.005 ;
        RECT 283.090 395.720 284.090 399.005 ;
        RECT 284.930 395.720 285.930 399.005 ;
        RECT 286.770 395.720 287.770 399.005 ;
        RECT 288.610 395.720 289.150 399.005 ;
        RECT 289.990 395.720 290.990 399.005 ;
        RECT 291.830 395.720 292.830 399.005 ;
        RECT 293.670 395.720 294.670 399.005 ;
        RECT 295.510 395.720 296.510 399.005 ;
        RECT 297.350 395.720 297.890 399.005 ;
        RECT 298.730 395.720 299.730 399.005 ;
        RECT 300.570 395.720 301.570 399.005 ;
        RECT 302.410 395.720 303.410 399.005 ;
        RECT 304.250 395.720 304.790 399.005 ;
        RECT 305.630 395.720 306.630 399.005 ;
        RECT 307.470 395.720 308.470 399.005 ;
        RECT 309.310 395.720 310.310 399.005 ;
        RECT 311.150 395.720 311.690 399.005 ;
        RECT 312.530 395.720 313.530 399.005 ;
        RECT 314.370 395.720 315.370 399.005 ;
        RECT 316.210 395.720 317.210 399.005 ;
        RECT 318.050 395.720 318.590 399.005 ;
        RECT 319.430 395.720 320.430 399.005 ;
        RECT 321.270 395.720 322.270 399.005 ;
        RECT 323.110 395.720 324.110 399.005 ;
        RECT 324.950 395.720 325.950 399.005 ;
        RECT 326.790 395.720 327.330 399.005 ;
        RECT 328.170 395.720 329.170 399.005 ;
        RECT 330.010 395.720 331.010 399.005 ;
        RECT 331.850 395.720 332.850 399.005 ;
        RECT 333.690 395.720 334.230 399.005 ;
        RECT 335.070 395.720 336.070 399.005 ;
        RECT 336.910 395.720 337.910 399.005 ;
        RECT 338.750 395.720 339.750 399.005 ;
        RECT 340.590 395.720 341.130 399.005 ;
        RECT 341.970 395.720 342.970 399.005 ;
        RECT 343.810 395.720 344.810 399.005 ;
        RECT 345.650 395.720 346.650 399.005 ;
        RECT 347.490 395.720 348.490 399.005 ;
        RECT 349.330 395.720 349.870 399.005 ;
        RECT 350.710 395.720 351.710 399.005 ;
        RECT 352.550 395.720 353.550 399.005 ;
        RECT 354.390 395.720 355.390 399.005 ;
        RECT 356.230 395.720 356.770 399.005 ;
        RECT 357.610 395.720 358.610 399.005 ;
        RECT 359.450 395.720 360.450 399.005 ;
        RECT 361.290 395.720 362.290 399.005 ;
        RECT 363.130 395.720 363.670 399.005 ;
        RECT 364.510 395.720 365.510 399.005 ;
        RECT 366.350 395.720 367.350 399.005 ;
        RECT 368.190 395.720 369.190 399.005 ;
        RECT 370.030 395.720 370.570 399.005 ;
        RECT 371.410 395.720 372.410 399.005 ;
        RECT 373.250 395.720 374.250 399.005 ;
        RECT 375.090 395.720 376.090 399.005 ;
        RECT 376.930 395.720 377.930 399.005 ;
        RECT 378.770 395.720 379.310 399.005 ;
        RECT 380.150 395.720 381.150 399.005 ;
        RECT 381.990 395.720 382.990 399.005 ;
        RECT 383.830 395.720 384.830 399.005 ;
        RECT 385.670 395.720 386.210 399.005 ;
        RECT 387.050 395.720 388.050 399.005 ;
        RECT 388.890 395.720 389.890 399.005 ;
        RECT 390.730 395.720 391.730 399.005 ;
        RECT 392.570 395.720 393.110 399.005 ;
        RECT 393.950 395.720 394.950 399.005 ;
        RECT 395.790 395.720 396.790 399.005 ;
        RECT 397.630 395.720 398.630 399.005 ;
        RECT 0.560 4.280 399.180 395.720 ;
        RECT 1.110 0.835 1.650 4.280 ;
        RECT 2.490 0.835 3.490 4.280 ;
        RECT 4.330 0.835 5.330 4.280 ;
        RECT 6.170 0.835 6.710 4.280 ;
        RECT 7.550 0.835 8.550 4.280 ;
        RECT 9.390 0.835 10.390 4.280 ;
        RECT 11.230 0.835 12.230 4.280 ;
        RECT 13.070 0.835 13.610 4.280 ;
        RECT 14.450 0.835 15.450 4.280 ;
        RECT 16.290 0.835 17.290 4.280 ;
        RECT 18.130 0.835 19.130 4.280 ;
        RECT 19.970 0.835 20.510 4.280 ;
        RECT 21.350 0.835 22.350 4.280 ;
        RECT 23.190 0.835 24.190 4.280 ;
        RECT 25.030 0.835 26.030 4.280 ;
        RECT 26.870 0.835 27.410 4.280 ;
        RECT 28.250 0.835 29.250 4.280 ;
        RECT 30.090 0.835 31.090 4.280 ;
        RECT 31.930 0.835 32.470 4.280 ;
        RECT 33.310 0.835 34.310 4.280 ;
        RECT 35.150 0.835 36.150 4.280 ;
        RECT 36.990 0.835 37.990 4.280 ;
        RECT 38.830 0.835 39.370 4.280 ;
        RECT 40.210 0.835 41.210 4.280 ;
        RECT 42.050 0.835 43.050 4.280 ;
        RECT 43.890 0.835 44.890 4.280 ;
        RECT 45.730 0.835 46.270 4.280 ;
        RECT 47.110 0.835 48.110 4.280 ;
        RECT 48.950 0.835 49.950 4.280 ;
        RECT 50.790 0.835 51.790 4.280 ;
        RECT 52.630 0.835 53.170 4.280 ;
        RECT 54.010 0.835 55.010 4.280 ;
        RECT 55.850 0.835 56.850 4.280 ;
        RECT 57.690 0.835 58.230 4.280 ;
        RECT 59.070 0.835 60.070 4.280 ;
        RECT 60.910 0.835 61.910 4.280 ;
        RECT 62.750 0.835 63.750 4.280 ;
        RECT 64.590 0.835 65.130 4.280 ;
        RECT 65.970 0.835 66.970 4.280 ;
        RECT 67.810 0.835 68.810 4.280 ;
        RECT 69.650 0.835 70.650 4.280 ;
        RECT 71.490 0.835 72.030 4.280 ;
        RECT 72.870 0.835 73.870 4.280 ;
        RECT 74.710 0.835 75.710 4.280 ;
        RECT 76.550 0.835 77.550 4.280 ;
        RECT 78.390 0.835 78.930 4.280 ;
        RECT 79.770 0.835 80.770 4.280 ;
        RECT 81.610 0.835 82.610 4.280 ;
        RECT 83.450 0.835 83.990 4.280 ;
        RECT 84.830 0.835 85.830 4.280 ;
        RECT 86.670 0.835 87.670 4.280 ;
        RECT 88.510 0.835 89.510 4.280 ;
        RECT 90.350 0.835 90.890 4.280 ;
        RECT 91.730 0.835 92.730 4.280 ;
        RECT 93.570 0.835 94.570 4.280 ;
        RECT 95.410 0.835 96.410 4.280 ;
        RECT 97.250 0.835 97.790 4.280 ;
        RECT 98.630 0.835 99.630 4.280 ;
        RECT 100.470 0.835 101.470 4.280 ;
        RECT 102.310 0.835 103.310 4.280 ;
        RECT 104.150 0.835 104.690 4.280 ;
        RECT 105.530 0.835 106.530 4.280 ;
        RECT 107.370 0.835 108.370 4.280 ;
        RECT 109.210 0.835 109.750 4.280 ;
        RECT 110.590 0.835 111.590 4.280 ;
        RECT 112.430 0.835 113.430 4.280 ;
        RECT 114.270 0.835 115.270 4.280 ;
        RECT 116.110 0.835 116.650 4.280 ;
        RECT 117.490 0.835 118.490 4.280 ;
        RECT 119.330 0.835 120.330 4.280 ;
        RECT 121.170 0.835 122.170 4.280 ;
        RECT 123.010 0.835 123.550 4.280 ;
        RECT 124.390 0.835 125.390 4.280 ;
        RECT 126.230 0.835 127.230 4.280 ;
        RECT 128.070 0.835 129.070 4.280 ;
        RECT 129.910 0.835 130.450 4.280 ;
        RECT 131.290 0.835 132.290 4.280 ;
        RECT 133.130 0.835 134.130 4.280 ;
        RECT 134.970 0.835 135.510 4.280 ;
        RECT 136.350 0.835 137.350 4.280 ;
        RECT 138.190 0.835 139.190 4.280 ;
        RECT 140.030 0.835 141.030 4.280 ;
        RECT 141.870 0.835 142.410 4.280 ;
        RECT 143.250 0.835 144.250 4.280 ;
        RECT 145.090 0.835 146.090 4.280 ;
        RECT 146.930 0.835 147.930 4.280 ;
        RECT 148.770 0.835 149.310 4.280 ;
        RECT 150.150 0.835 151.150 4.280 ;
        RECT 151.990 0.835 152.990 4.280 ;
        RECT 153.830 0.835 154.830 4.280 ;
        RECT 155.670 0.835 156.210 4.280 ;
        RECT 157.050 0.835 158.050 4.280 ;
        RECT 158.890 0.835 159.890 4.280 ;
        RECT 160.730 0.835 161.270 4.280 ;
        RECT 162.110 0.835 163.110 4.280 ;
        RECT 163.950 0.835 164.950 4.280 ;
        RECT 165.790 0.835 166.790 4.280 ;
        RECT 167.630 0.835 168.170 4.280 ;
        RECT 169.010 0.835 170.010 4.280 ;
        RECT 170.850 0.835 171.850 4.280 ;
        RECT 172.690 0.835 173.690 4.280 ;
        RECT 174.530 0.835 175.070 4.280 ;
        RECT 175.910 0.835 176.910 4.280 ;
        RECT 177.750 0.835 178.750 4.280 ;
        RECT 179.590 0.835 180.590 4.280 ;
        RECT 181.430 0.835 181.970 4.280 ;
        RECT 182.810 0.835 183.810 4.280 ;
        RECT 184.650 0.835 185.650 4.280 ;
        RECT 186.490 0.835 187.030 4.280 ;
        RECT 187.870 0.835 188.870 4.280 ;
        RECT 189.710 0.835 190.710 4.280 ;
        RECT 191.550 0.835 192.550 4.280 ;
        RECT 193.390 0.835 193.930 4.280 ;
        RECT 194.770 0.835 195.770 4.280 ;
        RECT 196.610 0.835 197.610 4.280 ;
        RECT 198.450 0.835 199.450 4.280 ;
        RECT 200.290 0.835 200.830 4.280 ;
        RECT 201.670 0.835 202.670 4.280 ;
        RECT 203.510 0.835 204.510 4.280 ;
        RECT 205.350 0.835 206.350 4.280 ;
        RECT 207.190 0.835 207.730 4.280 ;
        RECT 208.570 0.835 209.570 4.280 ;
        RECT 210.410 0.835 211.410 4.280 ;
        RECT 212.250 0.835 213.250 4.280 ;
        RECT 214.090 0.835 214.630 4.280 ;
        RECT 215.470 0.835 216.470 4.280 ;
        RECT 217.310 0.835 218.310 4.280 ;
        RECT 219.150 0.835 219.690 4.280 ;
        RECT 220.530 0.835 221.530 4.280 ;
        RECT 222.370 0.835 223.370 4.280 ;
        RECT 224.210 0.835 225.210 4.280 ;
        RECT 226.050 0.835 226.590 4.280 ;
        RECT 227.430 0.835 228.430 4.280 ;
        RECT 229.270 0.835 230.270 4.280 ;
        RECT 231.110 0.835 232.110 4.280 ;
        RECT 232.950 0.835 233.490 4.280 ;
        RECT 234.330 0.835 235.330 4.280 ;
        RECT 236.170 0.835 237.170 4.280 ;
        RECT 238.010 0.835 239.010 4.280 ;
        RECT 239.850 0.835 240.390 4.280 ;
        RECT 241.230 0.835 242.230 4.280 ;
        RECT 243.070 0.835 244.070 4.280 ;
        RECT 244.910 0.835 245.450 4.280 ;
        RECT 246.290 0.835 247.290 4.280 ;
        RECT 248.130 0.835 249.130 4.280 ;
        RECT 249.970 0.835 250.970 4.280 ;
        RECT 251.810 0.835 252.350 4.280 ;
        RECT 253.190 0.835 254.190 4.280 ;
        RECT 255.030 0.835 256.030 4.280 ;
        RECT 256.870 0.835 257.870 4.280 ;
        RECT 258.710 0.835 259.250 4.280 ;
        RECT 260.090 0.835 261.090 4.280 ;
        RECT 261.930 0.835 262.930 4.280 ;
        RECT 263.770 0.835 264.770 4.280 ;
        RECT 265.610 0.835 266.150 4.280 ;
        RECT 266.990 0.835 267.990 4.280 ;
        RECT 268.830 0.835 269.830 4.280 ;
        RECT 270.670 0.835 271.210 4.280 ;
        RECT 272.050 0.835 273.050 4.280 ;
        RECT 273.890 0.835 274.890 4.280 ;
        RECT 275.730 0.835 276.730 4.280 ;
        RECT 277.570 0.835 278.110 4.280 ;
        RECT 278.950 0.835 279.950 4.280 ;
        RECT 280.790 0.835 281.790 4.280 ;
        RECT 282.630 0.835 283.630 4.280 ;
        RECT 284.470 0.835 285.010 4.280 ;
        RECT 285.850 0.835 286.850 4.280 ;
        RECT 287.690 0.835 288.690 4.280 ;
        RECT 289.530 0.835 290.530 4.280 ;
        RECT 291.370 0.835 291.910 4.280 ;
        RECT 292.750 0.835 293.750 4.280 ;
        RECT 294.590 0.835 295.590 4.280 ;
        RECT 296.430 0.835 296.970 4.280 ;
        RECT 297.810 0.835 298.810 4.280 ;
        RECT 299.650 0.835 300.650 4.280 ;
        RECT 301.490 0.835 302.490 4.280 ;
        RECT 303.330 0.835 303.870 4.280 ;
        RECT 304.710 0.835 305.710 4.280 ;
        RECT 306.550 0.835 307.550 4.280 ;
        RECT 308.390 0.835 309.390 4.280 ;
        RECT 310.230 0.835 310.770 4.280 ;
        RECT 311.610 0.835 312.610 4.280 ;
        RECT 313.450 0.835 314.450 4.280 ;
        RECT 315.290 0.835 316.290 4.280 ;
        RECT 317.130 0.835 317.670 4.280 ;
        RECT 318.510 0.835 319.510 4.280 ;
        RECT 320.350 0.835 321.350 4.280 ;
        RECT 322.190 0.835 322.730 4.280 ;
        RECT 323.570 0.835 324.570 4.280 ;
        RECT 325.410 0.835 326.410 4.280 ;
        RECT 327.250 0.835 328.250 4.280 ;
        RECT 329.090 0.835 329.630 4.280 ;
        RECT 330.470 0.835 331.470 4.280 ;
        RECT 332.310 0.835 333.310 4.280 ;
        RECT 334.150 0.835 335.150 4.280 ;
        RECT 335.990 0.835 336.530 4.280 ;
        RECT 337.370 0.835 338.370 4.280 ;
        RECT 339.210 0.835 340.210 4.280 ;
        RECT 341.050 0.835 342.050 4.280 ;
        RECT 342.890 0.835 343.430 4.280 ;
        RECT 344.270 0.835 345.270 4.280 ;
        RECT 346.110 0.835 347.110 4.280 ;
        RECT 347.950 0.835 348.490 4.280 ;
        RECT 349.330 0.835 350.330 4.280 ;
        RECT 351.170 0.835 352.170 4.280 ;
        RECT 353.010 0.835 354.010 4.280 ;
        RECT 354.850 0.835 355.390 4.280 ;
        RECT 356.230 0.835 357.230 4.280 ;
        RECT 358.070 0.835 359.070 4.280 ;
        RECT 359.910 0.835 360.910 4.280 ;
        RECT 361.750 0.835 362.290 4.280 ;
        RECT 363.130 0.835 364.130 4.280 ;
        RECT 364.970 0.835 365.970 4.280 ;
        RECT 366.810 0.835 367.810 4.280 ;
        RECT 368.650 0.835 369.190 4.280 ;
        RECT 370.030 0.835 371.030 4.280 ;
        RECT 371.870 0.835 372.870 4.280 ;
        RECT 373.710 0.835 374.250 4.280 ;
        RECT 375.090 0.835 376.090 4.280 ;
        RECT 376.930 0.835 377.930 4.280 ;
        RECT 378.770 0.835 379.770 4.280 ;
        RECT 380.610 0.835 381.150 4.280 ;
        RECT 381.990 0.835 382.990 4.280 ;
        RECT 383.830 0.835 384.830 4.280 ;
        RECT 385.670 0.835 386.670 4.280 ;
        RECT 387.510 0.835 388.050 4.280 ;
        RECT 388.890 0.835 389.890 4.280 ;
        RECT 390.730 0.835 391.730 4.280 ;
        RECT 392.570 0.835 393.570 4.280 ;
        RECT 394.410 0.835 394.950 4.280 ;
        RECT 395.790 0.835 396.790 4.280 ;
        RECT 397.630 0.835 398.630 4.280 ;
      LAYER met3 ;
        RECT 4.400 398.120 395.600 398.985 ;
        RECT 4.000 397.480 395.600 398.120 ;
        RECT 4.400 396.760 395.600 397.480 ;
        RECT 4.400 396.120 396.000 396.760 ;
        RECT 4.400 394.720 395.600 396.120 ;
        RECT 4.000 394.080 395.600 394.720 ;
        RECT 4.400 392.000 395.600 394.080 ;
        RECT 4.400 391.360 396.000 392.000 ;
        RECT 4.400 391.320 395.600 391.360 ;
        RECT 4.000 390.680 395.600 391.320 ;
        RECT 4.400 388.600 395.600 390.680 ;
        RECT 4.400 387.960 396.000 388.600 ;
        RECT 4.400 387.920 395.600 387.960 ;
        RECT 4.000 387.280 395.600 387.920 ;
        RECT 4.400 384.520 395.600 387.280 ;
        RECT 4.000 383.880 395.600 384.520 ;
        RECT 4.400 383.840 395.600 383.880 ;
        RECT 4.400 383.200 396.000 383.840 ;
        RECT 4.400 381.120 395.600 383.200 ;
        RECT 4.000 380.480 395.600 381.120 ;
        RECT 4.400 379.080 395.600 380.480 ;
        RECT 4.000 378.440 396.000 379.080 ;
        RECT 4.400 375.680 395.600 378.440 ;
        RECT 4.000 375.040 396.000 375.680 ;
        RECT 4.400 372.280 395.600 375.040 ;
        RECT 4.000 371.640 395.600 372.280 ;
        RECT 4.400 370.920 395.600 371.640 ;
        RECT 4.400 370.280 396.000 370.920 ;
        RECT 4.400 368.880 395.600 370.280 ;
        RECT 4.000 368.240 395.600 368.880 ;
        RECT 4.400 366.160 395.600 368.240 ;
        RECT 4.400 365.520 396.000 366.160 ;
        RECT 4.400 365.480 395.600 365.520 ;
        RECT 4.000 364.840 395.600 365.480 ;
        RECT 4.400 362.760 395.600 364.840 ;
        RECT 4.400 362.120 396.000 362.760 ;
        RECT 4.400 362.080 395.600 362.120 ;
        RECT 4.000 361.440 395.600 362.080 ;
        RECT 4.400 360.040 395.600 361.440 ;
        RECT 4.000 359.400 395.600 360.040 ;
        RECT 4.400 358.000 395.600 359.400 ;
        RECT 4.400 357.360 396.000 358.000 ;
        RECT 4.400 356.640 395.600 357.360 ;
        RECT 4.000 356.000 395.600 356.640 ;
        RECT 4.400 354.600 395.600 356.000 ;
        RECT 4.400 353.960 396.000 354.600 ;
        RECT 4.400 353.240 395.600 353.960 ;
        RECT 4.000 352.600 395.600 353.240 ;
        RECT 4.400 349.840 395.600 352.600 ;
        RECT 4.000 349.200 396.000 349.840 ;
        RECT 4.400 346.440 395.600 349.200 ;
        RECT 4.000 345.800 395.600 346.440 ;
        RECT 4.400 345.080 395.600 345.800 ;
        RECT 4.400 344.440 396.000 345.080 ;
        RECT 4.400 343.040 395.600 344.440 ;
        RECT 4.000 342.400 395.600 343.040 ;
        RECT 4.400 341.680 395.600 342.400 ;
        RECT 4.400 341.040 396.000 341.680 ;
        RECT 4.400 341.000 395.600 341.040 ;
        RECT 4.000 340.360 395.600 341.000 ;
        RECT 4.400 337.600 395.600 340.360 ;
        RECT 4.000 336.960 395.600 337.600 ;
        RECT 4.400 336.920 395.600 336.960 ;
        RECT 4.400 336.280 396.000 336.920 ;
        RECT 4.400 334.200 395.600 336.280 ;
        RECT 4.000 333.560 395.600 334.200 ;
        RECT 4.400 332.160 395.600 333.560 ;
        RECT 4.400 331.520 396.000 332.160 ;
        RECT 4.400 330.800 395.600 331.520 ;
        RECT 4.000 330.160 395.600 330.800 ;
        RECT 4.400 328.760 395.600 330.160 ;
        RECT 4.400 328.120 396.000 328.760 ;
        RECT 4.400 327.400 395.600 328.120 ;
        RECT 4.000 326.760 395.600 327.400 ;
        RECT 4.400 324.000 395.600 326.760 ;
        RECT 4.000 323.360 396.000 324.000 ;
        RECT 4.400 321.960 395.600 323.360 ;
        RECT 4.000 321.320 395.600 321.960 ;
        RECT 4.400 320.600 395.600 321.320 ;
        RECT 4.400 319.960 396.000 320.600 ;
        RECT 4.400 318.560 395.600 319.960 ;
        RECT 4.000 317.920 395.600 318.560 ;
        RECT 4.400 315.840 395.600 317.920 ;
        RECT 4.400 315.200 396.000 315.840 ;
        RECT 4.400 315.160 395.600 315.200 ;
        RECT 4.000 314.520 395.600 315.160 ;
        RECT 4.400 311.760 395.600 314.520 ;
        RECT 4.000 311.120 395.600 311.760 ;
        RECT 4.400 311.080 395.600 311.120 ;
        RECT 4.400 310.440 396.000 311.080 ;
        RECT 4.400 308.360 395.600 310.440 ;
        RECT 4.000 307.720 395.600 308.360 ;
        RECT 4.400 307.680 395.600 307.720 ;
        RECT 4.400 307.040 396.000 307.680 ;
        RECT 4.400 304.960 395.600 307.040 ;
        RECT 4.000 304.320 395.600 304.960 ;
        RECT 4.400 302.920 395.600 304.320 ;
        RECT 4.000 302.280 396.000 302.920 ;
        RECT 4.400 299.520 395.600 302.280 ;
        RECT 4.000 298.880 395.600 299.520 ;
        RECT 4.400 298.160 395.600 298.880 ;
        RECT 4.400 297.520 396.000 298.160 ;
        RECT 4.400 296.120 395.600 297.520 ;
        RECT 4.000 295.480 395.600 296.120 ;
        RECT 4.400 294.760 395.600 295.480 ;
        RECT 4.400 294.120 396.000 294.760 ;
        RECT 4.400 292.720 395.600 294.120 ;
        RECT 4.000 292.080 395.600 292.720 ;
        RECT 4.400 290.000 395.600 292.080 ;
        RECT 4.400 289.360 396.000 290.000 ;
        RECT 4.400 289.320 395.600 289.360 ;
        RECT 4.000 288.680 395.600 289.320 ;
        RECT 4.400 286.600 395.600 288.680 ;
        RECT 4.400 285.960 396.000 286.600 ;
        RECT 4.400 285.920 395.600 285.960 ;
        RECT 4.000 285.280 395.600 285.920 ;
        RECT 4.400 283.880 395.600 285.280 ;
        RECT 4.000 283.240 395.600 283.880 ;
        RECT 4.400 281.840 395.600 283.240 ;
        RECT 4.400 281.200 396.000 281.840 ;
        RECT 4.400 280.480 395.600 281.200 ;
        RECT 4.000 279.840 395.600 280.480 ;
        RECT 4.400 277.080 395.600 279.840 ;
        RECT 4.000 276.440 396.000 277.080 ;
        RECT 4.400 273.680 395.600 276.440 ;
        RECT 4.000 273.040 396.000 273.680 ;
        RECT 4.400 270.280 395.600 273.040 ;
        RECT 4.000 269.640 395.600 270.280 ;
        RECT 4.400 268.920 395.600 269.640 ;
        RECT 4.400 268.280 396.000 268.920 ;
        RECT 4.400 266.880 395.600 268.280 ;
        RECT 4.000 266.240 395.600 266.880 ;
        RECT 4.400 264.840 395.600 266.240 ;
        RECT 4.000 264.200 395.600 264.840 ;
        RECT 4.400 264.160 395.600 264.200 ;
        RECT 4.400 263.520 396.000 264.160 ;
        RECT 4.400 261.440 395.600 263.520 ;
        RECT 4.000 260.800 395.600 261.440 ;
        RECT 4.400 260.760 395.600 260.800 ;
        RECT 4.400 260.120 396.000 260.760 ;
        RECT 4.400 258.040 395.600 260.120 ;
        RECT 4.000 257.400 395.600 258.040 ;
        RECT 4.400 256.000 395.600 257.400 ;
        RECT 4.400 255.360 396.000 256.000 ;
        RECT 4.400 254.640 395.600 255.360 ;
        RECT 4.000 254.000 395.600 254.640 ;
        RECT 4.400 252.600 395.600 254.000 ;
        RECT 4.400 251.960 396.000 252.600 ;
        RECT 4.400 251.240 395.600 251.960 ;
        RECT 4.000 250.600 395.600 251.240 ;
        RECT 4.400 247.840 395.600 250.600 ;
        RECT 4.000 247.200 396.000 247.840 ;
        RECT 4.400 245.800 395.600 247.200 ;
        RECT 4.000 245.160 395.600 245.800 ;
        RECT 4.400 243.080 395.600 245.160 ;
        RECT 4.400 242.440 396.000 243.080 ;
        RECT 4.400 242.400 395.600 242.440 ;
        RECT 4.000 241.760 395.600 242.400 ;
        RECT 4.400 239.680 395.600 241.760 ;
        RECT 4.400 239.040 396.000 239.680 ;
        RECT 4.400 239.000 395.600 239.040 ;
        RECT 4.000 238.360 395.600 239.000 ;
        RECT 4.400 235.600 395.600 238.360 ;
        RECT 4.000 234.960 395.600 235.600 ;
        RECT 4.400 234.920 395.600 234.960 ;
        RECT 4.400 234.280 396.000 234.920 ;
        RECT 4.400 232.200 395.600 234.280 ;
        RECT 4.000 231.560 395.600 232.200 ;
        RECT 4.400 230.160 395.600 231.560 ;
        RECT 4.400 229.520 396.000 230.160 ;
        RECT 4.400 228.800 395.600 229.520 ;
        RECT 4.000 228.160 395.600 228.800 ;
        RECT 4.400 226.760 395.600 228.160 ;
        RECT 4.000 226.120 396.000 226.760 ;
        RECT 4.400 223.360 395.600 226.120 ;
        RECT 4.000 222.720 395.600 223.360 ;
        RECT 4.400 222.000 395.600 222.720 ;
        RECT 4.400 221.360 396.000 222.000 ;
        RECT 4.400 219.960 395.600 221.360 ;
        RECT 4.000 219.320 395.600 219.960 ;
        RECT 4.400 218.600 395.600 219.320 ;
        RECT 4.400 217.960 396.000 218.600 ;
        RECT 4.400 216.560 395.600 217.960 ;
        RECT 4.000 215.920 395.600 216.560 ;
        RECT 4.400 213.840 395.600 215.920 ;
        RECT 4.400 213.200 396.000 213.840 ;
        RECT 4.400 213.160 395.600 213.200 ;
        RECT 4.000 212.520 395.600 213.160 ;
        RECT 4.400 209.760 395.600 212.520 ;
        RECT 4.000 209.120 395.600 209.760 ;
        RECT 4.400 209.080 395.600 209.120 ;
        RECT 4.400 208.440 396.000 209.080 ;
        RECT 4.400 207.720 395.600 208.440 ;
        RECT 4.000 207.080 395.600 207.720 ;
        RECT 4.400 205.680 395.600 207.080 ;
        RECT 4.400 205.040 396.000 205.680 ;
        RECT 4.400 204.320 395.600 205.040 ;
        RECT 4.000 203.680 395.600 204.320 ;
        RECT 4.400 200.920 395.600 203.680 ;
        RECT 4.000 200.280 396.000 200.920 ;
        RECT 4.400 197.520 395.600 200.280 ;
        RECT 4.000 196.880 395.600 197.520 ;
        RECT 4.400 196.160 395.600 196.880 ;
        RECT 4.400 195.520 396.000 196.160 ;
        RECT 4.400 194.120 395.600 195.520 ;
        RECT 4.000 193.480 395.600 194.120 ;
        RECT 4.400 192.760 395.600 193.480 ;
        RECT 4.400 192.120 396.000 192.760 ;
        RECT 4.400 190.720 395.600 192.120 ;
        RECT 4.000 190.080 395.600 190.720 ;
        RECT 4.400 188.680 395.600 190.080 ;
        RECT 4.000 188.040 395.600 188.680 ;
        RECT 4.400 188.000 395.600 188.040 ;
        RECT 4.400 187.360 396.000 188.000 ;
        RECT 4.400 185.280 395.600 187.360 ;
        RECT 4.000 184.640 395.600 185.280 ;
        RECT 4.400 183.240 395.600 184.640 ;
        RECT 4.400 182.600 396.000 183.240 ;
        RECT 4.400 181.880 395.600 182.600 ;
        RECT 4.000 181.240 395.600 181.880 ;
        RECT 4.400 179.840 395.600 181.240 ;
        RECT 4.400 179.200 396.000 179.840 ;
        RECT 4.400 178.480 395.600 179.200 ;
        RECT 4.000 177.840 395.600 178.480 ;
        RECT 4.400 175.080 395.600 177.840 ;
        RECT 4.000 174.440 396.000 175.080 ;
        RECT 4.400 171.680 395.600 174.440 ;
        RECT 4.000 171.040 396.000 171.680 ;
        RECT 4.400 169.640 395.600 171.040 ;
        RECT 4.000 169.000 395.600 169.640 ;
        RECT 4.400 166.920 395.600 169.000 ;
        RECT 4.400 166.280 396.000 166.920 ;
        RECT 4.400 166.240 395.600 166.280 ;
        RECT 4.000 165.600 395.600 166.240 ;
        RECT 4.400 162.840 395.600 165.600 ;
        RECT 4.000 162.200 395.600 162.840 ;
        RECT 4.400 162.160 395.600 162.200 ;
        RECT 4.400 161.520 396.000 162.160 ;
        RECT 4.400 159.440 395.600 161.520 ;
        RECT 4.000 158.800 395.600 159.440 ;
        RECT 4.400 158.760 395.600 158.800 ;
        RECT 4.400 158.120 396.000 158.760 ;
        RECT 4.400 156.040 395.600 158.120 ;
        RECT 4.000 155.400 395.600 156.040 ;
        RECT 4.400 154.000 395.600 155.400 ;
        RECT 4.400 153.360 396.000 154.000 ;
        RECT 4.400 152.640 395.600 153.360 ;
        RECT 4.000 152.000 395.600 152.640 ;
        RECT 4.400 150.600 395.600 152.000 ;
        RECT 4.000 149.960 395.600 150.600 ;
        RECT 4.400 149.240 395.600 149.960 ;
        RECT 4.400 148.600 396.000 149.240 ;
        RECT 4.400 147.200 395.600 148.600 ;
        RECT 4.000 146.560 395.600 147.200 ;
        RECT 4.400 145.840 395.600 146.560 ;
        RECT 4.400 145.200 396.000 145.840 ;
        RECT 4.400 143.800 395.600 145.200 ;
        RECT 4.000 143.160 395.600 143.800 ;
        RECT 4.400 141.080 395.600 143.160 ;
        RECT 4.400 140.440 396.000 141.080 ;
        RECT 4.400 140.400 395.600 140.440 ;
        RECT 4.000 139.760 395.600 140.400 ;
        RECT 4.400 137.680 395.600 139.760 ;
        RECT 4.400 137.040 396.000 137.680 ;
        RECT 4.400 137.000 395.600 137.040 ;
        RECT 4.000 136.360 395.600 137.000 ;
        RECT 4.400 133.600 395.600 136.360 ;
        RECT 4.000 132.960 395.600 133.600 ;
        RECT 4.400 132.920 395.600 132.960 ;
        RECT 4.400 132.280 396.000 132.920 ;
        RECT 4.400 131.560 395.600 132.280 ;
        RECT 4.000 130.920 395.600 131.560 ;
        RECT 4.400 128.160 395.600 130.920 ;
        RECT 4.000 127.520 396.000 128.160 ;
        RECT 4.400 124.760 395.600 127.520 ;
        RECT 4.000 124.120 396.000 124.760 ;
        RECT 4.400 121.360 395.600 124.120 ;
        RECT 4.000 120.720 395.600 121.360 ;
        RECT 4.400 120.000 395.600 120.720 ;
        RECT 4.400 119.360 396.000 120.000 ;
        RECT 4.400 117.960 395.600 119.360 ;
        RECT 4.000 117.320 395.600 117.960 ;
        RECT 4.400 115.240 395.600 117.320 ;
        RECT 4.400 114.600 396.000 115.240 ;
        RECT 4.400 114.560 395.600 114.600 ;
        RECT 4.000 113.920 395.600 114.560 ;
        RECT 4.400 112.520 395.600 113.920 ;
        RECT 4.000 111.880 395.600 112.520 ;
        RECT 4.400 111.840 395.600 111.880 ;
        RECT 4.400 111.200 396.000 111.840 ;
        RECT 4.400 109.120 395.600 111.200 ;
        RECT 4.000 108.480 395.600 109.120 ;
        RECT 4.400 107.080 395.600 108.480 ;
        RECT 4.400 106.440 396.000 107.080 ;
        RECT 4.400 105.720 395.600 106.440 ;
        RECT 4.000 105.080 395.600 105.720 ;
        RECT 4.400 103.680 395.600 105.080 ;
        RECT 4.400 103.040 396.000 103.680 ;
        RECT 4.400 102.320 395.600 103.040 ;
        RECT 4.000 101.680 395.600 102.320 ;
        RECT 4.400 98.920 395.600 101.680 ;
        RECT 4.000 98.280 396.000 98.920 ;
        RECT 4.400 95.520 395.600 98.280 ;
        RECT 4.000 94.880 395.600 95.520 ;
        RECT 4.400 94.160 395.600 94.880 ;
        RECT 4.400 93.520 396.000 94.160 ;
        RECT 4.400 93.480 395.600 93.520 ;
        RECT 4.000 92.840 395.600 93.480 ;
        RECT 4.400 90.760 395.600 92.840 ;
        RECT 4.400 90.120 396.000 90.760 ;
        RECT 4.400 90.080 395.600 90.120 ;
        RECT 4.000 89.440 395.600 90.080 ;
        RECT 4.400 86.680 395.600 89.440 ;
        RECT 4.000 86.040 395.600 86.680 ;
        RECT 4.400 86.000 395.600 86.040 ;
        RECT 4.400 85.360 396.000 86.000 ;
        RECT 4.400 83.280 395.600 85.360 ;
        RECT 4.000 82.640 395.600 83.280 ;
        RECT 4.400 81.240 395.600 82.640 ;
        RECT 4.400 80.600 396.000 81.240 ;
        RECT 4.400 79.880 395.600 80.600 ;
        RECT 4.000 79.240 395.600 79.880 ;
        RECT 4.400 77.840 395.600 79.240 ;
        RECT 4.400 77.200 396.000 77.840 ;
        RECT 4.400 76.480 395.600 77.200 ;
        RECT 4.000 75.840 395.600 76.480 ;
        RECT 4.400 74.440 395.600 75.840 ;
        RECT 4.000 73.800 395.600 74.440 ;
        RECT 4.400 73.080 395.600 73.800 ;
        RECT 4.400 72.440 396.000 73.080 ;
        RECT 4.400 71.040 395.600 72.440 ;
        RECT 4.000 70.400 395.600 71.040 ;
        RECT 4.400 69.680 395.600 70.400 ;
        RECT 4.400 69.040 396.000 69.680 ;
        RECT 4.400 67.640 395.600 69.040 ;
        RECT 4.000 67.000 395.600 67.640 ;
        RECT 4.400 64.920 395.600 67.000 ;
        RECT 4.400 64.280 396.000 64.920 ;
        RECT 4.400 64.240 395.600 64.280 ;
        RECT 4.000 63.600 395.600 64.240 ;
        RECT 4.400 60.840 395.600 63.600 ;
        RECT 4.000 60.200 395.600 60.840 ;
        RECT 4.400 60.160 395.600 60.200 ;
        RECT 4.400 59.520 396.000 60.160 ;
        RECT 4.400 57.440 395.600 59.520 ;
        RECT 4.000 56.800 395.600 57.440 ;
        RECT 4.400 56.760 395.600 56.800 ;
        RECT 4.400 56.120 396.000 56.760 ;
        RECT 4.400 55.400 395.600 56.120 ;
        RECT 4.000 54.760 395.600 55.400 ;
        RECT 4.400 52.000 395.600 54.760 ;
        RECT 4.000 51.360 396.000 52.000 ;
        RECT 4.400 48.600 395.600 51.360 ;
        RECT 4.000 47.960 395.600 48.600 ;
        RECT 4.400 47.240 395.600 47.960 ;
        RECT 4.400 46.600 396.000 47.240 ;
        RECT 4.400 45.200 395.600 46.600 ;
        RECT 4.000 44.560 395.600 45.200 ;
        RECT 4.400 43.840 395.600 44.560 ;
        RECT 4.400 43.200 396.000 43.840 ;
        RECT 4.400 41.800 395.600 43.200 ;
        RECT 4.000 41.160 395.600 41.800 ;
        RECT 4.400 39.080 395.600 41.160 ;
        RECT 4.400 38.440 396.000 39.080 ;
        RECT 4.400 38.400 395.600 38.440 ;
        RECT 4.000 37.760 395.600 38.400 ;
        RECT 4.400 36.360 395.600 37.760 ;
        RECT 4.000 35.720 395.600 36.360 ;
        RECT 4.400 35.680 395.600 35.720 ;
        RECT 4.400 35.040 396.000 35.680 ;
        RECT 4.400 32.960 395.600 35.040 ;
        RECT 4.000 32.320 395.600 32.960 ;
        RECT 4.400 30.920 395.600 32.320 ;
        RECT 4.400 30.280 396.000 30.920 ;
        RECT 4.400 29.560 395.600 30.280 ;
        RECT 4.000 28.920 395.600 29.560 ;
        RECT 4.400 26.160 395.600 28.920 ;
        RECT 4.000 25.520 396.000 26.160 ;
        RECT 4.400 22.760 395.600 25.520 ;
        RECT 4.000 22.120 396.000 22.760 ;
        RECT 4.400 19.360 395.600 22.120 ;
        RECT 4.000 18.720 395.600 19.360 ;
        RECT 4.400 18.000 395.600 18.720 ;
        RECT 4.400 17.360 396.000 18.000 ;
        RECT 4.400 17.320 395.600 17.360 ;
        RECT 4.000 16.680 395.600 17.320 ;
        RECT 4.400 13.920 395.600 16.680 ;
        RECT 4.000 13.280 395.600 13.920 ;
        RECT 4.400 13.240 395.600 13.280 ;
        RECT 4.400 12.600 396.000 13.240 ;
        RECT 4.400 10.520 395.600 12.600 ;
        RECT 4.000 9.880 395.600 10.520 ;
        RECT 4.400 9.840 395.600 9.880 ;
        RECT 4.400 9.200 396.000 9.840 ;
        RECT 4.400 7.120 395.600 9.200 ;
        RECT 4.000 6.480 395.600 7.120 ;
        RECT 4.400 5.080 395.600 6.480 ;
        RECT 4.400 4.440 396.000 5.080 ;
        RECT 4.400 3.720 395.600 4.440 ;
        RECT 4.000 3.080 395.600 3.720 ;
        RECT 4.400 0.855 395.600 3.080 ;
      LAYER met4 ;
        RECT 10.415 10.240 20.640 325.545 ;
        RECT 23.040 10.240 97.440 325.545 ;
        RECT 99.840 10.240 174.240 325.545 ;
        RECT 176.640 10.240 251.040 325.545 ;
        RECT 253.440 10.240 327.840 325.545 ;
        RECT 330.240 10.240 386.105 325.545 ;
        RECT 10.415 9.695 386.105 10.240 ;
  END
END chip_controller
END LIBRARY

