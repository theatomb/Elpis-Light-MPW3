VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 1496.000 9.110 1500.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.920 4.000 1286.520 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.770 1496.000 1292.050 1500.000 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.670 0.000 1298.950 4.000 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1263.480 1500.000 1264.080 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1317.880 4.000 1318.480 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1281.160 1500.000 1281.760 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1298.840 1500.000 1299.440 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1381.120 4.000 1381.720 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1315.840 1500.000 1316.440 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1396.760 4.000 1397.360 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1351.200 1500.000 1351.800 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.110 1496.000 1328.390 1500.000 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 1496.000 1346.330 1500.000 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.070 0.000 1386.350 4.000 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 1496.000 1364.270 1500.000 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1412.400 4.000 1413.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.040 4.000 1428.640 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.330 1496.000 1400.610 1500.000 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.510 0.000 1438.790 4.000 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1403.560 1500.000 1404.160 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1420.560 1500.000 1421.160 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1475.640 4.000 1476.240 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 1496.000 1436.490 1500.000 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.470 0.000 1473.750 4.000 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1455.920 1500.000 1456.520 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1490.600 1500.000 1491.200 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 1496.000 515.110 1500.000 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 287.000 1500.000 287.600 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 339.360 1500.000 339.960 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 25.200 1500.000 25.800 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 408.720 1500.000 409.320 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 1496.000 623.210 1500.000 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 548.800 1500.000 549.400 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 1496.000 713.830 1500.000 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 670.520 1500.000 671.120 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 1496.000 786.050 1500.000 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 705.880 1500.000 706.480 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 59.880 1500.000 60.480 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 740.560 1500.000 741.160 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 1496.000 822.390 1500.000 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.760 4.000 734.360 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 758.240 1500.000 758.840 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 1496.000 840.330 1500.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 775.240 1500.000 775.840 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 4.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 0.000 845.850 4.000 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.070 0.000 880.350 4.000 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 1496.000 948.890 1500.000 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 1496.000 966.830 1500.000 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 862.280 1500.000 862.880 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 77.560 1500.000 78.160 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 897.640 1500.000 898.240 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 914.640 1500.000 915.240 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 891.520 4.000 892.120 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.160 4.000 907.760 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 1496.000 1002.710 1500.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 967.000 1500.000 967.600 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1002.360 1500.000 1002.960 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 4.000 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 970.400 4.000 971.000 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 1496.000 262.110 1500.000 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 1496.000 1021.110 1500.000 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.770 1496.000 1039.050 1500.000 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1019.360 1500.000 1019.960 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1037.040 1500.000 1037.640 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1054.720 1500.000 1055.320 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.280 4.000 1049.880 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1071.720 1500.000 1072.320 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 1496.000 1093.330 1500.000 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 1496.000 297.990 1500.000 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 0.000 1072.630 4.000 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 1496.000 1147.610 1500.000 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1089.400 1500.000 1090.000 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 0.000 1107.130 4.000 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1112.520 4.000 1113.120 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1107.080 1500.000 1107.680 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1143.800 4.000 1144.400 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 1496.000 1183.490 1500.000 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1158.760 1500.000 1159.360 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1160.120 4.000 1160.720 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1496.000 315.930 1500.000 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 0.000 1124.610 4.000 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1176.440 1500.000 1177.040 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.810 0.000 1142.090 4.000 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1191.400 4.000 1192.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1194.120 1500.000 1194.720 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1211.120 1500.000 1211.720 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1223.360 4.000 1223.960 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.730 0.000 1212.010 4.000 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.210 0.000 1229.490 4.000 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 164.600 1500.000 165.200 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1496.000 135.610 1500.000 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 1496.000 424.490 1500.000 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 1496.000 478.770 1500.000 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 1496.000 496.710 1500.000 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 269.320 1500.000 269.920 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 304.680 1500.000 305.280 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 1496.000 568.930 1500.000 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 374.040 1500.000 374.640 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 426.400 1500.000 427.000 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 528.400 4.000 529.000 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 1496.000 641.610 1500.000 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 1496.000 659.550 1500.000 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 1496.000 677.490 1500.000 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 1496.000 695.430 1500.000 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 1496.000 171.490 1500.000 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 1496.000 768.110 1500.000 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 1496.000 207.830 1500.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 95.240 1500.000 95.840 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 1496.000 280.050 1500.000 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 147.600 1500.000 148.200 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 1496.000 334.330 1500.000 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 1496.000 81.330 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 1496.000 117.210 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 1496.000 99.270 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 182.280 1500.000 182.880 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 199.960 1500.000 200.560 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 357.040 1500.000 357.640 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 391.720 1500.000 392.320 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 42.880 1500.000 43.480 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 1496.000 243.710 1500.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 1496.000 352.270 1500.000 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 8.200 1500.000 8.800 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 0.000 1264.450 4.000 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1228.800 1500.000 1229.400 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 0.000 1281.930 4.000 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1246.480 1500.000 1247.080 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 0.000 1316.430 4.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1333.520 4.000 1334.120 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.160 4.000 1349.760 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1365.480 4.000 1366.080 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 0.000 1333.910 4.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1333.520 1500.000 1334.120 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 1496.000 1309.990 1500.000 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.110 0.000 1351.390 4.000 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1368.200 1500.000 1368.800 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.550 0.000 1403.830 4.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 1496.000 1382.210 1500.000 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 0.000 1421.310 4.000 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1444.360 4.000 1444.960 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1385.880 1500.000 1386.480 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 0.000 1456.270 4.000 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1496.000 460.830 1500.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1460.000 4.000 1460.600 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.270 1496.000 1418.550 1500.000 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.280 4.000 1491.880 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1438.240 1500.000 1438.840 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.610 1496.000 1454.890 1500.000 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.550 1496.000 1472.830 1500.000 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1472.920 1500.000 1473.520 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 1496.000 1490.770 1500.000 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 216.960 1500.000 217.560 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 234.640 1500.000 235.240 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 1496.000 533.050 1500.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 321.680 1500.000 322.280 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 444.080 1500.000 444.680 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 478.760 1500.000 479.360 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 513.440 1500.000 514.040 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 601.160 1500.000 601.760 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 1496.000 731.770 1500.000 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 635.840 1500.000 636.440 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 653.520 1500.000 654.120 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.880 4.000 655.480 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 1496.000 803.990 1500.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 688.200 1500.000 688.800 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 722.880 1500.000 723.480 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1496.000 225.770 1500.000 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 1496.000 858.270 1500.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 792.920 1500.000 793.520 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 1496.000 876.210 1500.000 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 0.000 793.410 4.000 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 4.000 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 1496.000 894.610 1500.000 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 809.920 1500.000 810.520 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 1496.000 912.550 1500.000 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 1496.000 930.490 1500.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.920 4.000 844.520 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 827.600 1500.000 828.200 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 845.280 1500.000 845.880 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 0.000 915.310 4.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 879.960 1500.000 880.560 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 0.000 932.790 4.000 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 1496.000 984.770 1500.000 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 932.320 1500.000 932.920 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.800 4.000 923.400 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 950.000 1500.000 950.600 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.760 4.000 955.360 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 984.680 1500.000 985.280 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 0.000 985.230 4.000 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 129.920 1500.000 130.520 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.680 4.000 1002.280 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 4.000 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.000 4.000 1018.600 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 1496.000 1056.990 1500.000 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 0.000 1020.190 4.000 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 1496.000 1075.390 1500.000 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 4.000 1065.520 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.870 0.000 1055.150 4.000 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 1496.000 1111.270 1500.000 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930 1496.000 1129.210 1500.000 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 0.000 1089.650 4.000 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.270 1496.000 1165.550 1500.000 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.880 4.000 1097.480 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.160 4.000 1128.760 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1124.080 1500.000 1124.680 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1141.760 1500.000 1142.360 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.610 1496.000 1201.890 1500.000 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 1496.000 1219.830 1500.000 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.490 1496.000 1237.770 1500.000 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 1496.000 370.210 1500.000 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.430 1496.000 1255.710 1500.000 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1175.760 4.000 1176.360 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.040 4.000 1207.640 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 4.000 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 1496.000 1274.110 1500.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.000 4.000 1239.600 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.280 4.000 1270.880 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 0.000 1246.970 4.000 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 1496.000 388.610 1500.000 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 1496.000 44.990 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 1496.000 62.930 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 1496.000 153.550 1500.000 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 1496.000 442.430 1500.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 252.320 1500.000 252.920 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1496.000 550.990 1500.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 1496.000 587.330 1500.000 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 1496.000 605.270 1500.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 461.080 1500.000 461.680 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 496.440 1500.000 497.040 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 531.120 1500.000 531.720 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 565.800 1500.000 566.400 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 583.480 1500.000 584.080 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 618.160 1500.000 618.760 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 1496.000 189.430 1500.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 1496.000 749.710 1500.000 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 112.240 1500.000 112.840 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 1496.000 406.550 1500.000 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 1496.000 27.050 1500.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.080 1488.080 ;
      LAYER met2 ;
        RECT 6.990 1495.720 8.550 1496.410 ;
        RECT 9.390 1495.720 26.490 1496.410 ;
        RECT 27.330 1495.720 44.430 1496.410 ;
        RECT 45.270 1495.720 62.370 1496.410 ;
        RECT 63.210 1495.720 80.770 1496.410 ;
        RECT 81.610 1495.720 98.710 1496.410 ;
        RECT 99.550 1495.720 116.650 1496.410 ;
        RECT 117.490 1495.720 135.050 1496.410 ;
        RECT 135.890 1495.720 152.990 1496.410 ;
        RECT 153.830 1495.720 170.930 1496.410 ;
        RECT 171.770 1495.720 188.870 1496.410 ;
        RECT 189.710 1495.720 207.270 1496.410 ;
        RECT 208.110 1495.720 225.210 1496.410 ;
        RECT 226.050 1495.720 243.150 1496.410 ;
        RECT 243.990 1495.720 261.550 1496.410 ;
        RECT 262.390 1495.720 279.490 1496.410 ;
        RECT 280.330 1495.720 297.430 1496.410 ;
        RECT 298.270 1495.720 315.370 1496.410 ;
        RECT 316.210 1495.720 333.770 1496.410 ;
        RECT 334.610 1495.720 351.710 1496.410 ;
        RECT 352.550 1495.720 369.650 1496.410 ;
        RECT 370.490 1495.720 388.050 1496.410 ;
        RECT 388.890 1495.720 405.990 1496.410 ;
        RECT 406.830 1495.720 423.930 1496.410 ;
        RECT 424.770 1495.720 441.870 1496.410 ;
        RECT 442.710 1495.720 460.270 1496.410 ;
        RECT 461.110 1495.720 478.210 1496.410 ;
        RECT 479.050 1495.720 496.150 1496.410 ;
        RECT 496.990 1495.720 514.550 1496.410 ;
        RECT 515.390 1495.720 532.490 1496.410 ;
        RECT 533.330 1495.720 550.430 1496.410 ;
        RECT 551.270 1495.720 568.370 1496.410 ;
        RECT 569.210 1495.720 586.770 1496.410 ;
        RECT 587.610 1495.720 604.710 1496.410 ;
        RECT 605.550 1495.720 622.650 1496.410 ;
        RECT 623.490 1495.720 641.050 1496.410 ;
        RECT 641.890 1495.720 658.990 1496.410 ;
        RECT 659.830 1495.720 676.930 1496.410 ;
        RECT 677.770 1495.720 694.870 1496.410 ;
        RECT 695.710 1495.720 713.270 1496.410 ;
        RECT 714.110 1495.720 731.210 1496.410 ;
        RECT 732.050 1495.720 749.150 1496.410 ;
        RECT 749.990 1495.720 767.550 1496.410 ;
        RECT 768.390 1495.720 785.490 1496.410 ;
        RECT 786.330 1495.720 803.430 1496.410 ;
        RECT 804.270 1495.720 821.830 1496.410 ;
        RECT 822.670 1495.720 839.770 1496.410 ;
        RECT 840.610 1495.720 857.710 1496.410 ;
        RECT 858.550 1495.720 875.650 1496.410 ;
        RECT 876.490 1495.720 894.050 1496.410 ;
        RECT 894.890 1495.720 911.990 1496.410 ;
        RECT 912.830 1495.720 929.930 1496.410 ;
        RECT 930.770 1495.720 948.330 1496.410 ;
        RECT 949.170 1495.720 966.270 1496.410 ;
        RECT 967.110 1495.720 984.210 1496.410 ;
        RECT 985.050 1495.720 1002.150 1496.410 ;
        RECT 1002.990 1495.720 1020.550 1496.410 ;
        RECT 1021.390 1495.720 1038.490 1496.410 ;
        RECT 1039.330 1495.720 1056.430 1496.410 ;
        RECT 1057.270 1495.720 1074.830 1496.410 ;
        RECT 1075.670 1495.720 1092.770 1496.410 ;
        RECT 1093.610 1495.720 1110.710 1496.410 ;
        RECT 1111.550 1495.720 1128.650 1496.410 ;
        RECT 1129.490 1495.720 1147.050 1496.410 ;
        RECT 1147.890 1495.720 1164.990 1496.410 ;
        RECT 1165.830 1495.720 1182.930 1496.410 ;
        RECT 1183.770 1495.720 1201.330 1496.410 ;
        RECT 1202.170 1495.720 1219.270 1496.410 ;
        RECT 1220.110 1495.720 1237.210 1496.410 ;
        RECT 1238.050 1495.720 1255.150 1496.410 ;
        RECT 1255.990 1495.720 1273.550 1496.410 ;
        RECT 1274.390 1495.720 1291.490 1496.410 ;
        RECT 1292.330 1495.720 1309.430 1496.410 ;
        RECT 1310.270 1495.720 1327.830 1496.410 ;
        RECT 1328.670 1495.720 1345.770 1496.410 ;
        RECT 1346.610 1495.720 1363.710 1496.410 ;
        RECT 1364.550 1495.720 1381.650 1496.410 ;
        RECT 1382.490 1495.720 1400.050 1496.410 ;
        RECT 1400.890 1495.720 1417.990 1496.410 ;
        RECT 1418.830 1495.720 1435.930 1496.410 ;
        RECT 1436.770 1495.720 1454.330 1496.410 ;
        RECT 1455.170 1495.720 1472.270 1496.410 ;
        RECT 1473.110 1495.720 1490.210 1496.410 ;
        RECT 1491.050 1495.720 1491.220 1496.410 ;
        RECT 6.990 4.280 1491.220 1495.720 ;
        RECT 6.990 4.000 8.090 4.280 ;
        RECT 8.930 4.000 25.110 4.280 ;
        RECT 25.950 4.000 42.590 4.280 ;
        RECT 43.430 4.000 60.070 4.280 ;
        RECT 60.910 4.000 77.550 4.280 ;
        RECT 78.390 4.000 95.030 4.280 ;
        RECT 95.870 4.000 112.510 4.280 ;
        RECT 113.350 4.000 129.990 4.280 ;
        RECT 130.830 4.000 147.470 4.280 ;
        RECT 148.310 4.000 164.950 4.280 ;
        RECT 165.790 4.000 182.430 4.280 ;
        RECT 183.270 4.000 199.910 4.280 ;
        RECT 200.750 4.000 217.390 4.280 ;
        RECT 218.230 4.000 234.410 4.280 ;
        RECT 235.250 4.000 251.890 4.280 ;
        RECT 252.730 4.000 269.370 4.280 ;
        RECT 270.210 4.000 286.850 4.280 ;
        RECT 287.690 4.000 304.330 4.280 ;
        RECT 305.170 4.000 321.810 4.280 ;
        RECT 322.650 4.000 339.290 4.280 ;
        RECT 340.130 4.000 356.770 4.280 ;
        RECT 357.610 4.000 374.250 4.280 ;
        RECT 375.090 4.000 391.730 4.280 ;
        RECT 392.570 4.000 409.210 4.280 ;
        RECT 410.050 4.000 426.690 4.280 ;
        RECT 427.530 4.000 443.710 4.280 ;
        RECT 444.550 4.000 461.190 4.280 ;
        RECT 462.030 4.000 478.670 4.280 ;
        RECT 479.510 4.000 496.150 4.280 ;
        RECT 496.990 4.000 513.630 4.280 ;
        RECT 514.470 4.000 531.110 4.280 ;
        RECT 531.950 4.000 548.590 4.280 ;
        RECT 549.430 4.000 566.070 4.280 ;
        RECT 566.910 4.000 583.550 4.280 ;
        RECT 584.390 4.000 601.030 4.280 ;
        RECT 601.870 4.000 618.510 4.280 ;
        RECT 619.350 4.000 635.990 4.280 ;
        RECT 636.830 4.000 653.010 4.280 ;
        RECT 653.850 4.000 670.490 4.280 ;
        RECT 671.330 4.000 687.970 4.280 ;
        RECT 688.810 4.000 705.450 4.280 ;
        RECT 706.290 4.000 722.930 4.280 ;
        RECT 723.770 4.000 740.410 4.280 ;
        RECT 741.250 4.000 757.890 4.280 ;
        RECT 758.730 4.000 775.370 4.280 ;
        RECT 776.210 4.000 792.850 4.280 ;
        RECT 793.690 4.000 810.330 4.280 ;
        RECT 811.170 4.000 827.810 4.280 ;
        RECT 828.650 4.000 845.290 4.280 ;
        RECT 846.130 4.000 862.770 4.280 ;
        RECT 863.610 4.000 879.790 4.280 ;
        RECT 880.630 4.000 897.270 4.280 ;
        RECT 898.110 4.000 914.750 4.280 ;
        RECT 915.590 4.000 932.230 4.280 ;
        RECT 933.070 4.000 949.710 4.280 ;
        RECT 950.550 4.000 967.190 4.280 ;
        RECT 968.030 4.000 984.670 4.280 ;
        RECT 985.510 4.000 1002.150 4.280 ;
        RECT 1002.990 4.000 1019.630 4.280 ;
        RECT 1020.470 4.000 1037.110 4.280 ;
        RECT 1037.950 4.000 1054.590 4.280 ;
        RECT 1055.430 4.000 1072.070 4.280 ;
        RECT 1072.910 4.000 1089.090 4.280 ;
        RECT 1089.930 4.000 1106.570 4.280 ;
        RECT 1107.410 4.000 1124.050 4.280 ;
        RECT 1124.890 4.000 1141.530 4.280 ;
        RECT 1142.370 4.000 1159.010 4.280 ;
        RECT 1159.850 4.000 1176.490 4.280 ;
        RECT 1177.330 4.000 1193.970 4.280 ;
        RECT 1194.810 4.000 1211.450 4.280 ;
        RECT 1212.290 4.000 1228.930 4.280 ;
        RECT 1229.770 4.000 1246.410 4.280 ;
        RECT 1247.250 4.000 1263.890 4.280 ;
        RECT 1264.730 4.000 1281.370 4.280 ;
        RECT 1282.210 4.000 1298.390 4.280 ;
        RECT 1299.230 4.000 1315.870 4.280 ;
        RECT 1316.710 4.000 1333.350 4.280 ;
        RECT 1334.190 4.000 1350.830 4.280 ;
        RECT 1351.670 4.000 1368.310 4.280 ;
        RECT 1369.150 4.000 1385.790 4.280 ;
        RECT 1386.630 4.000 1403.270 4.280 ;
        RECT 1404.110 4.000 1420.750 4.280 ;
        RECT 1421.590 4.000 1438.230 4.280 ;
        RECT 1439.070 4.000 1455.710 4.280 ;
        RECT 1456.550 4.000 1473.190 4.280 ;
        RECT 1474.030 4.000 1490.670 4.280 ;
      LAYER met3 ;
        RECT 4.400 1491.600 1496.000 1491.745 ;
        RECT 4.400 1490.880 1495.600 1491.600 ;
        RECT 4.000 1490.200 1495.600 1490.880 ;
        RECT 4.000 1476.640 1496.000 1490.200 ;
        RECT 4.400 1475.240 1496.000 1476.640 ;
        RECT 4.000 1473.920 1496.000 1475.240 ;
        RECT 4.000 1472.520 1495.600 1473.920 ;
        RECT 4.000 1461.000 1496.000 1472.520 ;
        RECT 4.400 1459.600 1496.000 1461.000 ;
        RECT 4.000 1456.920 1496.000 1459.600 ;
        RECT 4.000 1455.520 1495.600 1456.920 ;
        RECT 4.000 1445.360 1496.000 1455.520 ;
        RECT 4.400 1443.960 1496.000 1445.360 ;
        RECT 4.000 1439.240 1496.000 1443.960 ;
        RECT 4.000 1437.840 1495.600 1439.240 ;
        RECT 4.000 1429.040 1496.000 1437.840 ;
        RECT 4.400 1427.640 1496.000 1429.040 ;
        RECT 4.000 1421.560 1496.000 1427.640 ;
        RECT 4.000 1420.160 1495.600 1421.560 ;
        RECT 4.000 1413.400 1496.000 1420.160 ;
        RECT 4.400 1412.000 1496.000 1413.400 ;
        RECT 4.000 1404.560 1496.000 1412.000 ;
        RECT 4.000 1403.160 1495.600 1404.560 ;
        RECT 4.000 1397.760 1496.000 1403.160 ;
        RECT 4.400 1396.360 1496.000 1397.760 ;
        RECT 4.000 1386.880 1496.000 1396.360 ;
        RECT 4.000 1385.480 1495.600 1386.880 ;
        RECT 4.000 1382.120 1496.000 1385.480 ;
        RECT 4.400 1380.720 1496.000 1382.120 ;
        RECT 4.000 1369.200 1496.000 1380.720 ;
        RECT 4.000 1367.800 1495.600 1369.200 ;
        RECT 4.000 1366.480 1496.000 1367.800 ;
        RECT 4.400 1365.080 1496.000 1366.480 ;
        RECT 4.000 1352.200 1496.000 1365.080 ;
        RECT 4.000 1350.800 1495.600 1352.200 ;
        RECT 4.000 1350.160 1496.000 1350.800 ;
        RECT 4.400 1348.760 1496.000 1350.160 ;
        RECT 4.000 1334.520 1496.000 1348.760 ;
        RECT 4.400 1333.120 1495.600 1334.520 ;
        RECT 4.000 1318.880 1496.000 1333.120 ;
        RECT 4.400 1317.480 1496.000 1318.880 ;
        RECT 4.000 1316.840 1496.000 1317.480 ;
        RECT 4.000 1315.440 1495.600 1316.840 ;
        RECT 4.000 1303.240 1496.000 1315.440 ;
        RECT 4.400 1301.840 1496.000 1303.240 ;
        RECT 4.000 1299.840 1496.000 1301.840 ;
        RECT 4.000 1298.440 1495.600 1299.840 ;
        RECT 4.000 1286.920 1496.000 1298.440 ;
        RECT 4.400 1285.520 1496.000 1286.920 ;
        RECT 4.000 1282.160 1496.000 1285.520 ;
        RECT 4.000 1280.760 1495.600 1282.160 ;
        RECT 4.000 1271.280 1496.000 1280.760 ;
        RECT 4.400 1269.880 1496.000 1271.280 ;
        RECT 4.000 1264.480 1496.000 1269.880 ;
        RECT 4.000 1263.080 1495.600 1264.480 ;
        RECT 4.000 1255.640 1496.000 1263.080 ;
        RECT 4.400 1254.240 1496.000 1255.640 ;
        RECT 4.000 1247.480 1496.000 1254.240 ;
        RECT 4.000 1246.080 1495.600 1247.480 ;
        RECT 4.000 1240.000 1496.000 1246.080 ;
        RECT 4.400 1238.600 1496.000 1240.000 ;
        RECT 4.000 1229.800 1496.000 1238.600 ;
        RECT 4.000 1228.400 1495.600 1229.800 ;
        RECT 4.000 1224.360 1496.000 1228.400 ;
        RECT 4.400 1222.960 1496.000 1224.360 ;
        RECT 4.000 1212.120 1496.000 1222.960 ;
        RECT 4.000 1210.720 1495.600 1212.120 ;
        RECT 4.000 1208.040 1496.000 1210.720 ;
        RECT 4.400 1206.640 1496.000 1208.040 ;
        RECT 4.000 1195.120 1496.000 1206.640 ;
        RECT 4.000 1193.720 1495.600 1195.120 ;
        RECT 4.000 1192.400 1496.000 1193.720 ;
        RECT 4.400 1191.000 1496.000 1192.400 ;
        RECT 4.000 1177.440 1496.000 1191.000 ;
        RECT 4.000 1176.760 1495.600 1177.440 ;
        RECT 4.400 1176.040 1495.600 1176.760 ;
        RECT 4.400 1175.360 1496.000 1176.040 ;
        RECT 4.000 1161.120 1496.000 1175.360 ;
        RECT 4.400 1159.760 1496.000 1161.120 ;
        RECT 4.400 1159.720 1495.600 1159.760 ;
        RECT 4.000 1158.360 1495.600 1159.720 ;
        RECT 4.000 1144.800 1496.000 1158.360 ;
        RECT 4.400 1143.400 1496.000 1144.800 ;
        RECT 4.000 1142.760 1496.000 1143.400 ;
        RECT 4.000 1141.360 1495.600 1142.760 ;
        RECT 4.000 1129.160 1496.000 1141.360 ;
        RECT 4.400 1127.760 1496.000 1129.160 ;
        RECT 4.000 1125.080 1496.000 1127.760 ;
        RECT 4.000 1123.680 1495.600 1125.080 ;
        RECT 4.000 1113.520 1496.000 1123.680 ;
        RECT 4.400 1112.120 1496.000 1113.520 ;
        RECT 4.000 1108.080 1496.000 1112.120 ;
        RECT 4.000 1106.680 1495.600 1108.080 ;
        RECT 4.000 1097.880 1496.000 1106.680 ;
        RECT 4.400 1096.480 1496.000 1097.880 ;
        RECT 4.000 1090.400 1496.000 1096.480 ;
        RECT 4.000 1089.000 1495.600 1090.400 ;
        RECT 4.000 1082.240 1496.000 1089.000 ;
        RECT 4.400 1080.840 1496.000 1082.240 ;
        RECT 4.000 1072.720 1496.000 1080.840 ;
        RECT 4.000 1071.320 1495.600 1072.720 ;
        RECT 4.000 1065.920 1496.000 1071.320 ;
        RECT 4.400 1064.520 1496.000 1065.920 ;
        RECT 4.000 1055.720 1496.000 1064.520 ;
        RECT 4.000 1054.320 1495.600 1055.720 ;
        RECT 4.000 1050.280 1496.000 1054.320 ;
        RECT 4.400 1048.880 1496.000 1050.280 ;
        RECT 4.000 1038.040 1496.000 1048.880 ;
        RECT 4.000 1036.640 1495.600 1038.040 ;
        RECT 4.000 1034.640 1496.000 1036.640 ;
        RECT 4.400 1033.240 1496.000 1034.640 ;
        RECT 4.000 1020.360 1496.000 1033.240 ;
        RECT 4.000 1019.000 1495.600 1020.360 ;
        RECT 4.400 1018.960 1495.600 1019.000 ;
        RECT 4.400 1017.600 1496.000 1018.960 ;
        RECT 4.000 1003.360 1496.000 1017.600 ;
        RECT 4.000 1002.680 1495.600 1003.360 ;
        RECT 4.400 1001.960 1495.600 1002.680 ;
        RECT 4.400 1001.280 1496.000 1001.960 ;
        RECT 4.000 987.040 1496.000 1001.280 ;
        RECT 4.400 985.680 1496.000 987.040 ;
        RECT 4.400 985.640 1495.600 985.680 ;
        RECT 4.000 984.280 1495.600 985.640 ;
        RECT 4.000 971.400 1496.000 984.280 ;
        RECT 4.400 970.000 1496.000 971.400 ;
        RECT 4.000 968.000 1496.000 970.000 ;
        RECT 4.000 966.600 1495.600 968.000 ;
        RECT 4.000 955.760 1496.000 966.600 ;
        RECT 4.400 954.360 1496.000 955.760 ;
        RECT 4.000 951.000 1496.000 954.360 ;
        RECT 4.000 949.600 1495.600 951.000 ;
        RECT 4.000 940.120 1496.000 949.600 ;
        RECT 4.400 938.720 1496.000 940.120 ;
        RECT 4.000 933.320 1496.000 938.720 ;
        RECT 4.000 931.920 1495.600 933.320 ;
        RECT 4.000 923.800 1496.000 931.920 ;
        RECT 4.400 922.400 1496.000 923.800 ;
        RECT 4.000 915.640 1496.000 922.400 ;
        RECT 4.000 914.240 1495.600 915.640 ;
        RECT 4.000 908.160 1496.000 914.240 ;
        RECT 4.400 906.760 1496.000 908.160 ;
        RECT 4.000 898.640 1496.000 906.760 ;
        RECT 4.000 897.240 1495.600 898.640 ;
        RECT 4.000 892.520 1496.000 897.240 ;
        RECT 4.400 891.120 1496.000 892.520 ;
        RECT 4.000 880.960 1496.000 891.120 ;
        RECT 4.000 879.560 1495.600 880.960 ;
        RECT 4.000 876.880 1496.000 879.560 ;
        RECT 4.400 875.480 1496.000 876.880 ;
        RECT 4.000 863.280 1496.000 875.480 ;
        RECT 4.000 861.880 1495.600 863.280 ;
        RECT 4.000 860.560 1496.000 861.880 ;
        RECT 4.400 859.160 1496.000 860.560 ;
        RECT 4.000 846.280 1496.000 859.160 ;
        RECT 4.000 844.920 1495.600 846.280 ;
        RECT 4.400 844.880 1495.600 844.920 ;
        RECT 4.400 843.520 1496.000 844.880 ;
        RECT 4.000 829.280 1496.000 843.520 ;
        RECT 4.400 828.600 1496.000 829.280 ;
        RECT 4.400 827.880 1495.600 828.600 ;
        RECT 4.000 827.200 1495.600 827.880 ;
        RECT 4.000 813.640 1496.000 827.200 ;
        RECT 4.400 812.240 1496.000 813.640 ;
        RECT 4.000 810.920 1496.000 812.240 ;
        RECT 4.000 809.520 1495.600 810.920 ;
        RECT 4.000 798.000 1496.000 809.520 ;
        RECT 4.400 796.600 1496.000 798.000 ;
        RECT 4.000 793.920 1496.000 796.600 ;
        RECT 4.000 792.520 1495.600 793.920 ;
        RECT 4.000 781.680 1496.000 792.520 ;
        RECT 4.400 780.280 1496.000 781.680 ;
        RECT 4.000 776.240 1496.000 780.280 ;
        RECT 4.000 774.840 1495.600 776.240 ;
        RECT 4.000 766.040 1496.000 774.840 ;
        RECT 4.400 764.640 1496.000 766.040 ;
        RECT 4.000 759.240 1496.000 764.640 ;
        RECT 4.000 757.840 1495.600 759.240 ;
        RECT 4.000 750.400 1496.000 757.840 ;
        RECT 4.400 749.000 1496.000 750.400 ;
        RECT 4.000 741.560 1496.000 749.000 ;
        RECT 4.000 740.160 1495.600 741.560 ;
        RECT 4.000 734.760 1496.000 740.160 ;
        RECT 4.400 733.360 1496.000 734.760 ;
        RECT 4.000 723.880 1496.000 733.360 ;
        RECT 4.000 722.480 1495.600 723.880 ;
        RECT 4.000 718.440 1496.000 722.480 ;
        RECT 4.400 717.040 1496.000 718.440 ;
        RECT 4.000 706.880 1496.000 717.040 ;
        RECT 4.000 705.480 1495.600 706.880 ;
        RECT 4.000 702.800 1496.000 705.480 ;
        RECT 4.400 701.400 1496.000 702.800 ;
        RECT 4.000 689.200 1496.000 701.400 ;
        RECT 4.000 687.800 1495.600 689.200 ;
        RECT 4.000 687.160 1496.000 687.800 ;
        RECT 4.400 685.760 1496.000 687.160 ;
        RECT 4.000 671.520 1496.000 685.760 ;
        RECT 4.400 670.120 1495.600 671.520 ;
        RECT 4.000 655.880 1496.000 670.120 ;
        RECT 4.400 654.520 1496.000 655.880 ;
        RECT 4.400 654.480 1495.600 654.520 ;
        RECT 4.000 653.120 1495.600 654.480 ;
        RECT 4.000 639.560 1496.000 653.120 ;
        RECT 4.400 638.160 1496.000 639.560 ;
        RECT 4.000 636.840 1496.000 638.160 ;
        RECT 4.000 635.440 1495.600 636.840 ;
        RECT 4.000 623.920 1496.000 635.440 ;
        RECT 4.400 622.520 1496.000 623.920 ;
        RECT 4.000 619.160 1496.000 622.520 ;
        RECT 4.000 617.760 1495.600 619.160 ;
        RECT 4.000 608.280 1496.000 617.760 ;
        RECT 4.400 606.880 1496.000 608.280 ;
        RECT 4.000 602.160 1496.000 606.880 ;
        RECT 4.000 600.760 1495.600 602.160 ;
        RECT 4.000 592.640 1496.000 600.760 ;
        RECT 4.400 591.240 1496.000 592.640 ;
        RECT 4.000 584.480 1496.000 591.240 ;
        RECT 4.000 583.080 1495.600 584.480 ;
        RECT 4.000 576.320 1496.000 583.080 ;
        RECT 4.400 574.920 1496.000 576.320 ;
        RECT 4.000 566.800 1496.000 574.920 ;
        RECT 4.000 565.400 1495.600 566.800 ;
        RECT 4.000 560.680 1496.000 565.400 ;
        RECT 4.400 559.280 1496.000 560.680 ;
        RECT 4.000 549.800 1496.000 559.280 ;
        RECT 4.000 548.400 1495.600 549.800 ;
        RECT 4.000 545.040 1496.000 548.400 ;
        RECT 4.400 543.640 1496.000 545.040 ;
        RECT 4.000 532.120 1496.000 543.640 ;
        RECT 4.000 530.720 1495.600 532.120 ;
        RECT 4.000 529.400 1496.000 530.720 ;
        RECT 4.400 528.000 1496.000 529.400 ;
        RECT 4.000 514.440 1496.000 528.000 ;
        RECT 4.000 513.760 1495.600 514.440 ;
        RECT 4.400 513.040 1495.600 513.760 ;
        RECT 4.400 512.360 1496.000 513.040 ;
        RECT 4.000 497.440 1496.000 512.360 ;
        RECT 4.400 496.040 1495.600 497.440 ;
        RECT 4.000 481.800 1496.000 496.040 ;
        RECT 4.400 480.400 1496.000 481.800 ;
        RECT 4.000 479.760 1496.000 480.400 ;
        RECT 4.000 478.360 1495.600 479.760 ;
        RECT 4.000 466.160 1496.000 478.360 ;
        RECT 4.400 464.760 1496.000 466.160 ;
        RECT 4.000 462.080 1496.000 464.760 ;
        RECT 4.000 460.680 1495.600 462.080 ;
        RECT 4.000 450.520 1496.000 460.680 ;
        RECT 4.400 449.120 1496.000 450.520 ;
        RECT 4.000 445.080 1496.000 449.120 ;
        RECT 4.000 443.680 1495.600 445.080 ;
        RECT 4.000 434.200 1496.000 443.680 ;
        RECT 4.400 432.800 1496.000 434.200 ;
        RECT 4.000 427.400 1496.000 432.800 ;
        RECT 4.000 426.000 1495.600 427.400 ;
        RECT 4.000 418.560 1496.000 426.000 ;
        RECT 4.400 417.160 1496.000 418.560 ;
        RECT 4.000 409.720 1496.000 417.160 ;
        RECT 4.000 408.320 1495.600 409.720 ;
        RECT 4.000 402.920 1496.000 408.320 ;
        RECT 4.400 401.520 1496.000 402.920 ;
        RECT 4.000 392.720 1496.000 401.520 ;
        RECT 4.000 391.320 1495.600 392.720 ;
        RECT 4.000 387.280 1496.000 391.320 ;
        RECT 4.400 385.880 1496.000 387.280 ;
        RECT 4.000 375.040 1496.000 385.880 ;
        RECT 4.000 373.640 1495.600 375.040 ;
        RECT 4.000 371.640 1496.000 373.640 ;
        RECT 4.400 370.240 1496.000 371.640 ;
        RECT 4.000 358.040 1496.000 370.240 ;
        RECT 4.000 356.640 1495.600 358.040 ;
        RECT 4.000 355.320 1496.000 356.640 ;
        RECT 4.400 353.920 1496.000 355.320 ;
        RECT 4.000 340.360 1496.000 353.920 ;
        RECT 4.000 339.680 1495.600 340.360 ;
        RECT 4.400 338.960 1495.600 339.680 ;
        RECT 4.400 338.280 1496.000 338.960 ;
        RECT 4.000 324.040 1496.000 338.280 ;
        RECT 4.400 322.680 1496.000 324.040 ;
        RECT 4.400 322.640 1495.600 322.680 ;
        RECT 4.000 321.280 1495.600 322.640 ;
        RECT 4.000 308.400 1496.000 321.280 ;
        RECT 4.400 307.000 1496.000 308.400 ;
        RECT 4.000 305.680 1496.000 307.000 ;
        RECT 4.000 304.280 1495.600 305.680 ;
        RECT 4.000 292.080 1496.000 304.280 ;
        RECT 4.400 290.680 1496.000 292.080 ;
        RECT 4.000 288.000 1496.000 290.680 ;
        RECT 4.000 286.600 1495.600 288.000 ;
        RECT 4.000 276.440 1496.000 286.600 ;
        RECT 4.400 275.040 1496.000 276.440 ;
        RECT 4.000 270.320 1496.000 275.040 ;
        RECT 4.000 268.920 1495.600 270.320 ;
        RECT 4.000 260.800 1496.000 268.920 ;
        RECT 4.400 259.400 1496.000 260.800 ;
        RECT 4.000 253.320 1496.000 259.400 ;
        RECT 4.000 251.920 1495.600 253.320 ;
        RECT 4.000 245.160 1496.000 251.920 ;
        RECT 4.400 243.760 1496.000 245.160 ;
        RECT 4.000 235.640 1496.000 243.760 ;
        RECT 4.000 234.240 1495.600 235.640 ;
        RECT 4.000 229.520 1496.000 234.240 ;
        RECT 4.400 228.120 1496.000 229.520 ;
        RECT 4.000 217.960 1496.000 228.120 ;
        RECT 4.000 216.560 1495.600 217.960 ;
        RECT 4.000 213.200 1496.000 216.560 ;
        RECT 4.400 211.800 1496.000 213.200 ;
        RECT 4.000 200.960 1496.000 211.800 ;
        RECT 4.000 199.560 1495.600 200.960 ;
        RECT 4.000 197.560 1496.000 199.560 ;
        RECT 4.400 196.160 1496.000 197.560 ;
        RECT 4.000 183.280 1496.000 196.160 ;
        RECT 4.000 181.920 1495.600 183.280 ;
        RECT 4.400 181.880 1495.600 181.920 ;
        RECT 4.400 180.520 1496.000 181.880 ;
        RECT 4.000 166.280 1496.000 180.520 ;
        RECT 4.400 165.600 1496.000 166.280 ;
        RECT 4.400 164.880 1495.600 165.600 ;
        RECT 4.000 164.200 1495.600 164.880 ;
        RECT 4.000 149.960 1496.000 164.200 ;
        RECT 4.400 148.600 1496.000 149.960 ;
        RECT 4.400 148.560 1495.600 148.600 ;
        RECT 4.000 147.200 1495.600 148.560 ;
        RECT 4.000 134.320 1496.000 147.200 ;
        RECT 4.400 132.920 1496.000 134.320 ;
        RECT 4.000 130.920 1496.000 132.920 ;
        RECT 4.000 129.520 1495.600 130.920 ;
        RECT 4.000 118.680 1496.000 129.520 ;
        RECT 4.400 117.280 1496.000 118.680 ;
        RECT 4.000 113.240 1496.000 117.280 ;
        RECT 4.000 111.840 1495.600 113.240 ;
        RECT 4.000 103.040 1496.000 111.840 ;
        RECT 4.400 101.640 1496.000 103.040 ;
        RECT 4.000 96.240 1496.000 101.640 ;
        RECT 4.000 94.840 1495.600 96.240 ;
        RECT 4.000 87.400 1496.000 94.840 ;
        RECT 4.400 86.000 1496.000 87.400 ;
        RECT 4.000 78.560 1496.000 86.000 ;
        RECT 4.000 77.160 1495.600 78.560 ;
        RECT 4.000 71.080 1496.000 77.160 ;
        RECT 4.400 69.680 1496.000 71.080 ;
        RECT 4.000 60.880 1496.000 69.680 ;
        RECT 4.000 59.480 1495.600 60.880 ;
        RECT 4.000 55.440 1496.000 59.480 ;
        RECT 4.400 54.040 1496.000 55.440 ;
        RECT 4.000 43.880 1496.000 54.040 ;
        RECT 4.000 42.480 1495.600 43.880 ;
        RECT 4.000 39.800 1496.000 42.480 ;
        RECT 4.400 38.400 1496.000 39.800 ;
        RECT 4.000 26.200 1496.000 38.400 ;
        RECT 4.000 24.800 1495.600 26.200 ;
        RECT 4.000 24.160 1496.000 24.800 ;
        RECT 4.400 22.760 1496.000 24.160 ;
        RECT 4.000 9.200 1496.000 22.760 ;
        RECT 4.000 8.520 1495.600 9.200 ;
        RECT 4.400 7.800 1495.600 8.520 ;
        RECT 4.400 7.655 1496.000 7.800 ;
      LAYER met4 ;
        RECT 96.895 17.855 97.440 1485.625 ;
        RECT 99.840 17.855 174.240 1485.625 ;
        RECT 176.640 17.855 251.040 1485.625 ;
        RECT 253.440 17.855 327.840 1485.625 ;
        RECT 330.240 17.855 404.640 1485.625 ;
        RECT 407.040 17.855 481.440 1485.625 ;
        RECT 483.840 17.855 558.240 1485.625 ;
        RECT 560.640 17.855 635.040 1485.625 ;
        RECT 637.440 17.855 711.840 1485.625 ;
        RECT 714.240 17.855 788.640 1485.625 ;
        RECT 791.040 17.855 865.440 1485.625 ;
        RECT 867.840 17.855 942.240 1485.625 ;
        RECT 944.640 17.855 1019.040 1485.625 ;
        RECT 1021.440 17.855 1073.345 1485.625 ;
  END
END core
END LIBRARY

