VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1496.000 6.810 1500.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.840 4.000 1265.440 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 1496.000 1314.130 1500.000 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1283.880 4.000 1284.480 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1239.000 1500.000 1239.600 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 1496.000 1341.270 1500.000 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 0.000 1289.290 4.000 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.790 1496.000 1355.070 1500.000 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 1496.000 1368.870 1500.000 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.590 0.000 1322.870 4.000 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1280.480 1500.000 1281.080 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 1496.000 295.690 1500.000 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1301.560 1500.000 1302.160 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1322.640 1500.000 1323.240 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1358.680 4.000 1359.280 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1343.040 1500.000 1343.640 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1364.120 1500.000 1364.720 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 0.000 1407.510 4.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.790 1496.000 1424.070 1500.000 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.790 0.000 1424.070 4.000 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1405.600 1500.000 1406.200 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 1496.000 350.430 1500.000 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.390 1496.000 1451.670 1500.000 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1426.680 1500.000 1427.280 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1433.480 4.000 1434.080 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1468.160 1500.000 1468.760 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1457.830 0.000 1458.110 4.000 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.390 0.000 1474.670 4.000 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1470.880 4.000 1471.480 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 1496.000 1493.070 1500.000 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 426.400 1500.000 427.000 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 1496.000 433.230 1500.000 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 488.960 1500.000 489.560 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 1496.000 502.230 1500.000 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 1496.000 144.350 1500.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 635.160 1500.000 635.760 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 1496.000 529.370 1500.000 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 1496.000 584.570 1500.000 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 1496.000 653.570 1500.000 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 780.680 1500.000 781.280 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 1496.000 722.110 1500.000 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 1496.000 749.710 1500.000 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 702.480 4.000 703.080 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 1496.000 777.310 1500.000 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 93.200 1500.000 93.800 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 843.240 1500.000 843.840 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 1496.000 804.910 1500.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 1496.000 818.710 1500.000 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.280 4.000 777.880 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 796.320 4.000 796.920 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 864.320 1500.000 864.920 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 1496.000 845.850 1500.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 1496.000 226.690 1500.000 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 884.720 1500.000 885.320 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 1496.000 873.450 1500.000 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 1496.000 901.050 1500.000 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 1496.000 914.850 1500.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 926.880 1500.000 927.480 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.720 4.000 834.320 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.120 4.000 871.720 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.370 1496.000 928.650 1500.000 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 1496.000 942.450 1500.000 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 1496.000 956.250 1500.000 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 0.000 918.530 4.000 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 1496.000 983.850 1500.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.370 1496.000 997.650 1500.000 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 0.000 969.130 4.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 4.000 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.710 1496.000 1010.990 1500.000 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 1496.000 1038.590 1500.000 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 968.360 1500.000 968.960 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1021.400 4.000 1022.000 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.470 0.000 1036.750 4.000 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 0.000 1053.310 4.000 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 989.440 1500.000 990.040 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1058.800 4.000 1059.400 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1009.840 1500.000 1010.440 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.050 0.000 1070.330 4.000 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.200 4.000 1096.800 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.310 1496.000 1107.590 1500.000 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1051.320 1500.000 1051.920 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1114.560 4.000 1115.160 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1093.480 1500.000 1094.080 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 1496.000 1162.790 1500.000 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1113.880 1500.000 1114.480 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 1496.000 1176.130 1500.000 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1156.040 1500.000 1156.640 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.230 0.000 1154.510 4.000 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 239.400 1500.000 240.000 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1496.000 1217.530 1500.000 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.250 0.000 1171.530 4.000 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.650 1496.000 1258.930 1500.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1171.000 4.000 1171.600 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.830 0.000 1205.110 4.000 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.050 1496.000 1300.330 1500.000 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1245.800 4.000 1246.400 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1197.520 1500.000 1198.120 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 322.360 1500.000 322.960 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 1496.000 130.550 1500.000 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 1496.000 309.490 1500.000 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 384.920 1500.000 385.520 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1496.000 364.230 1500.000 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 447.480 1500.000 448.080 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1496.000 460.830 1500.000 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 1496.000 488.430 1500.000 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 530.440 1500.000 531.040 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 1496.000 158.150 1500.000 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 593.000 1500.000 593.600 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.760 4.000 496.360 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 676.640 1500.000 677.240 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 697.720 1500.000 698.320 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 1496.000 625.970 1500.000 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 1496.000 667.370 1500.000 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 1496.000 694.510 1500.000 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 1496.000 185.290 1500.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 134.680 1500.000 135.280 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 176.840 1500.000 177.440 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 259.800 1500.000 260.400 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1496.000 61.550 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 1496.000 102.950 1500.000 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 1496.000 89.150 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 1496.000 116.750 1500.000 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 1496.000 75.350 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 10.240 1500.000 10.840 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 1496.000 323.290 1500.000 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 1496.000 391.830 1500.000 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 468.560 1500.000 469.160 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 114.280 1500.000 114.880 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 1496.000 254.290 1500.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 1496.000 268.090 1500.000 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 280.880 1500.000 281.480 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 343.440 1500.000 344.040 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.410 0.000 1238.690 4.000 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.430 0.000 1255.710 4.000 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.650 1496.000 1327.930 1500.000 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 0.000 1272.730 4.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1321.280 4.000 1321.880 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1339.640 4.000 1340.240 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.030 0.000 1306.310 4.000 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1260.080 1500.000 1260.680 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1339.610 0.000 1339.890 4.000 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.630 0.000 1356.910 4.000 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.190 0.000 1373.470 4.000 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.210 0.000 1390.490 4.000 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.390 1496.000 1382.670 1500.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.190 1496.000 1396.470 1500.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.990 1496.000 1410.270 1500.000 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1385.200 1500.000 1385.800 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.590 1496.000 1437.870 1500.000 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1396.080 4.000 1396.680 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.810 0.000 1441.090 4.000 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1415.120 4.000 1415.720 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1447.760 1500.000 1448.360 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 1496.000 1465.470 1500.000 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1489.240 1500.000 1489.840 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1452.520 4.000 1453.120 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.990 1496.000 1479.270 1500.000 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.920 4.000 1490.520 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 0.000 1491.690 4.000 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 1496.000 405.630 1500.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 1496.000 447.030 1500.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 1496.000 474.630 1500.000 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 510.040 1500.000 510.640 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 551.520 1500.000 552.120 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 51.720 1500.000 52.320 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 655.560 1500.000 656.160 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 1496.000 598.370 1500.000 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 718.120 1500.000 718.720 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 4.000 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 739.200 1500.000 739.800 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 1496.000 708.310 1500.000 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 801.760 1500.000 802.360 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 1496.000 735.910 1500.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1496.000 763.510 1500.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 1496.000 791.110 1500.000 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 1496.000 199.090 1500.000 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 822.160 1500.000 822.760 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 0.000 716.130 4.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.230 1496.000 832.510 1500.000 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 1496.000 240.490 1500.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.370 1496.000 859.650 1500.000 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 1496.000 887.250 1500.000 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 905.800 1500.000 906.400 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 0.000 800.770 4.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.080 4.000 852.680 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.160 4.000 890.760 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 908.520 4.000 909.120 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 0.000 884.950 4.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 927.560 4.000 928.160 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.920 4.000 946.520 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 1496.000 970.050 1500.000 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.270 0.000 935.550 4.000 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.830 0.000 952.110 4.000 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.870 0.000 986.150 4.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 947.280 1500.000 947.880 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.510 1496.000 1024.790 1500.000 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 1496.000 1052.390 1500.000 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 1496.000 281.890 1500.000 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.960 4.000 965.560 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1002.360 4.000 1002.960 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.450 0.000 1019.730 4.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1039.760 4.000 1040.360 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 1496.000 1066.190 1500.000 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 1496.000 1079.990 1500.000 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.160 4.000 1077.760 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.510 1496.000 1093.790 1500.000 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.610 0.000 1086.890 4.000 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1030.920 1500.000 1031.520 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 197.240 1500.000 197.840 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 1496.000 1121.390 1500.000 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1072.400 1500.000 1073.000 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 1496.000 1135.190 1500.000 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.710 1496.000 1148.990 1500.000 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1133.600 4.000 1134.200 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.630 0.000 1103.910 4.000 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.650 1496.000 1189.930 1500.000 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1134.960 1500.000 1135.560 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 4.000 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.450 1496.000 1203.730 1500.000 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 301.280 1500.000 301.880 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 1496.000 1231.330 1500.000 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.850 1496.000 1245.130 1500.000 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 0.000 1188.090 4.000 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 1496.000 1272.730 1500.000 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1208.400 4.000 1209.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.250 1496.000 1286.530 1500.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1176.440 1500.000 1177.040 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.850 0.000 1222.130 4.000 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1218.600 1500.000 1219.200 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 363.840 1500.000 364.440 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 1496.000 33.950 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 1496.000 47.750 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 30.640 1500.000 31.240 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 1496.000 337.090 1500.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 406.000 1500.000 406.600 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 1496.000 378.030 1500.000 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 1496.000 419.430 1500.000 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.960 4.000 421.560 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 72.120 1500.000 72.720 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 572.600 1500.000 573.200 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 614.080 1500.000 614.680 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 1496.000 515.570 1500.000 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 1496.000 543.170 1500.000 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 1496.000 556.970 1500.000 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 1496.000 570.770 1500.000 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1496.000 612.170 1500.000 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 1496.000 639.770 1500.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 1496.000 171.950 1500.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 1496.000 680.710 1500.000 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 760.280 1500.000 760.880 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1496.000 212.890 1500.000 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 155.760 1500.000 156.360 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 218.320 1500.000 218.920 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 1496.000 20.150 1500.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.080 1488.820 ;
      LAYER met2 ;
        RECT 7.090 1495.720 19.590 1496.410 ;
        RECT 20.430 1495.720 33.390 1496.410 ;
        RECT 34.230 1495.720 47.190 1496.410 ;
        RECT 48.030 1495.720 60.990 1496.410 ;
        RECT 61.830 1495.720 74.790 1496.410 ;
        RECT 75.630 1495.720 88.590 1496.410 ;
        RECT 89.430 1495.720 102.390 1496.410 ;
        RECT 103.230 1495.720 116.190 1496.410 ;
        RECT 117.030 1495.720 129.990 1496.410 ;
        RECT 130.830 1495.720 143.790 1496.410 ;
        RECT 144.630 1495.720 157.590 1496.410 ;
        RECT 158.430 1495.720 171.390 1496.410 ;
        RECT 172.230 1495.720 184.730 1496.410 ;
        RECT 185.570 1495.720 198.530 1496.410 ;
        RECT 199.370 1495.720 212.330 1496.410 ;
        RECT 213.170 1495.720 226.130 1496.410 ;
        RECT 226.970 1495.720 239.930 1496.410 ;
        RECT 240.770 1495.720 253.730 1496.410 ;
        RECT 254.570 1495.720 267.530 1496.410 ;
        RECT 268.370 1495.720 281.330 1496.410 ;
        RECT 282.170 1495.720 295.130 1496.410 ;
        RECT 295.970 1495.720 308.930 1496.410 ;
        RECT 309.770 1495.720 322.730 1496.410 ;
        RECT 323.570 1495.720 336.530 1496.410 ;
        RECT 337.370 1495.720 349.870 1496.410 ;
        RECT 350.710 1495.720 363.670 1496.410 ;
        RECT 364.510 1495.720 377.470 1496.410 ;
        RECT 378.310 1495.720 391.270 1496.410 ;
        RECT 392.110 1495.720 405.070 1496.410 ;
        RECT 405.910 1495.720 418.870 1496.410 ;
        RECT 419.710 1495.720 432.670 1496.410 ;
        RECT 433.510 1495.720 446.470 1496.410 ;
        RECT 447.310 1495.720 460.270 1496.410 ;
        RECT 461.110 1495.720 474.070 1496.410 ;
        RECT 474.910 1495.720 487.870 1496.410 ;
        RECT 488.710 1495.720 501.670 1496.410 ;
        RECT 502.510 1495.720 515.010 1496.410 ;
        RECT 515.850 1495.720 528.810 1496.410 ;
        RECT 529.650 1495.720 542.610 1496.410 ;
        RECT 543.450 1495.720 556.410 1496.410 ;
        RECT 557.250 1495.720 570.210 1496.410 ;
        RECT 571.050 1495.720 584.010 1496.410 ;
        RECT 584.850 1495.720 597.810 1496.410 ;
        RECT 598.650 1495.720 611.610 1496.410 ;
        RECT 612.450 1495.720 625.410 1496.410 ;
        RECT 626.250 1495.720 639.210 1496.410 ;
        RECT 640.050 1495.720 653.010 1496.410 ;
        RECT 653.850 1495.720 666.810 1496.410 ;
        RECT 667.650 1495.720 680.150 1496.410 ;
        RECT 680.990 1495.720 693.950 1496.410 ;
        RECT 694.790 1495.720 707.750 1496.410 ;
        RECT 708.590 1495.720 721.550 1496.410 ;
        RECT 722.390 1495.720 735.350 1496.410 ;
        RECT 736.190 1495.720 749.150 1496.410 ;
        RECT 749.990 1495.720 762.950 1496.410 ;
        RECT 763.790 1495.720 776.750 1496.410 ;
        RECT 777.590 1495.720 790.550 1496.410 ;
        RECT 791.390 1495.720 804.350 1496.410 ;
        RECT 805.190 1495.720 818.150 1496.410 ;
        RECT 818.990 1495.720 831.950 1496.410 ;
        RECT 832.790 1495.720 845.290 1496.410 ;
        RECT 846.130 1495.720 859.090 1496.410 ;
        RECT 859.930 1495.720 872.890 1496.410 ;
        RECT 873.730 1495.720 886.690 1496.410 ;
        RECT 887.530 1495.720 900.490 1496.410 ;
        RECT 901.330 1495.720 914.290 1496.410 ;
        RECT 915.130 1495.720 928.090 1496.410 ;
        RECT 928.930 1495.720 941.890 1496.410 ;
        RECT 942.730 1495.720 955.690 1496.410 ;
        RECT 956.530 1495.720 969.490 1496.410 ;
        RECT 970.330 1495.720 983.290 1496.410 ;
        RECT 984.130 1495.720 997.090 1496.410 ;
        RECT 997.930 1495.720 1010.430 1496.410 ;
        RECT 1011.270 1495.720 1024.230 1496.410 ;
        RECT 1025.070 1495.720 1038.030 1496.410 ;
        RECT 1038.870 1495.720 1051.830 1496.410 ;
        RECT 1052.670 1495.720 1065.630 1496.410 ;
        RECT 1066.470 1495.720 1079.430 1496.410 ;
        RECT 1080.270 1495.720 1093.230 1496.410 ;
        RECT 1094.070 1495.720 1107.030 1496.410 ;
        RECT 1107.870 1495.720 1120.830 1496.410 ;
        RECT 1121.670 1495.720 1134.630 1496.410 ;
        RECT 1135.470 1495.720 1148.430 1496.410 ;
        RECT 1149.270 1495.720 1162.230 1496.410 ;
        RECT 1163.070 1495.720 1175.570 1496.410 ;
        RECT 1176.410 1495.720 1189.370 1496.410 ;
        RECT 1190.210 1495.720 1203.170 1496.410 ;
        RECT 1204.010 1495.720 1216.970 1496.410 ;
        RECT 1217.810 1495.720 1230.770 1496.410 ;
        RECT 1231.610 1495.720 1244.570 1496.410 ;
        RECT 1245.410 1495.720 1258.370 1496.410 ;
        RECT 1259.210 1495.720 1272.170 1496.410 ;
        RECT 1273.010 1495.720 1285.970 1496.410 ;
        RECT 1286.810 1495.720 1299.770 1496.410 ;
        RECT 1300.610 1495.720 1313.570 1496.410 ;
        RECT 1314.410 1495.720 1327.370 1496.410 ;
        RECT 1328.210 1495.720 1340.710 1496.410 ;
        RECT 1341.550 1495.720 1354.510 1496.410 ;
        RECT 1355.350 1495.720 1368.310 1496.410 ;
        RECT 1369.150 1495.720 1382.110 1496.410 ;
        RECT 1382.950 1495.720 1395.910 1496.410 ;
        RECT 1396.750 1495.720 1409.710 1496.410 ;
        RECT 1410.550 1495.720 1423.510 1496.410 ;
        RECT 1424.350 1495.720 1437.310 1496.410 ;
        RECT 1438.150 1495.720 1451.110 1496.410 ;
        RECT 1451.950 1495.720 1464.910 1496.410 ;
        RECT 1465.750 1495.720 1478.710 1496.410 ;
        RECT 1479.550 1495.720 1492.510 1496.410 ;
        RECT 6.540 4.280 1493.060 1495.720 ;
        RECT 6.540 3.670 8.090 4.280 ;
        RECT 8.930 3.670 24.650 4.280 ;
        RECT 25.490 3.670 41.670 4.280 ;
        RECT 42.510 3.670 58.230 4.280 ;
        RECT 59.070 3.670 75.250 4.280 ;
        RECT 76.090 3.670 92.270 4.280 ;
        RECT 93.110 3.670 108.830 4.280 ;
        RECT 109.670 3.670 125.850 4.280 ;
        RECT 126.690 3.670 142.870 4.280 ;
        RECT 143.710 3.670 159.430 4.280 ;
        RECT 160.270 3.670 176.450 4.280 ;
        RECT 177.290 3.670 193.470 4.280 ;
        RECT 194.310 3.670 210.030 4.280 ;
        RECT 210.870 3.670 227.050 4.280 ;
        RECT 227.890 3.670 243.610 4.280 ;
        RECT 244.450 3.670 260.630 4.280 ;
        RECT 261.470 3.670 277.650 4.280 ;
        RECT 278.490 3.670 294.210 4.280 ;
        RECT 295.050 3.670 311.230 4.280 ;
        RECT 312.070 3.670 328.250 4.280 ;
        RECT 329.090 3.670 344.810 4.280 ;
        RECT 345.650 3.670 361.830 4.280 ;
        RECT 362.670 3.670 378.850 4.280 ;
        RECT 379.690 3.670 395.410 4.280 ;
        RECT 396.250 3.670 412.430 4.280 ;
        RECT 413.270 3.670 429.450 4.280 ;
        RECT 430.290 3.670 446.010 4.280 ;
        RECT 446.850 3.670 463.030 4.280 ;
        RECT 463.870 3.670 479.590 4.280 ;
        RECT 480.430 3.670 496.610 4.280 ;
        RECT 497.450 3.670 513.630 4.280 ;
        RECT 514.470 3.670 530.190 4.280 ;
        RECT 531.030 3.670 547.210 4.280 ;
        RECT 548.050 3.670 564.230 4.280 ;
        RECT 565.070 3.670 580.790 4.280 ;
        RECT 581.630 3.670 597.810 4.280 ;
        RECT 598.650 3.670 614.830 4.280 ;
        RECT 615.670 3.670 631.390 4.280 ;
        RECT 632.230 3.670 648.410 4.280 ;
        RECT 649.250 3.670 664.970 4.280 ;
        RECT 665.810 3.670 681.990 4.280 ;
        RECT 682.830 3.670 699.010 4.280 ;
        RECT 699.850 3.670 715.570 4.280 ;
        RECT 716.410 3.670 732.590 4.280 ;
        RECT 733.430 3.670 749.610 4.280 ;
        RECT 750.450 3.670 766.170 4.280 ;
        RECT 767.010 3.670 783.190 4.280 ;
        RECT 784.030 3.670 800.210 4.280 ;
        RECT 801.050 3.670 816.770 4.280 ;
        RECT 817.610 3.670 833.790 4.280 ;
        RECT 834.630 3.670 850.810 4.280 ;
        RECT 851.650 3.670 867.370 4.280 ;
        RECT 868.210 3.670 884.390 4.280 ;
        RECT 885.230 3.670 900.950 4.280 ;
        RECT 901.790 3.670 917.970 4.280 ;
        RECT 918.810 3.670 934.990 4.280 ;
        RECT 935.830 3.670 951.550 4.280 ;
        RECT 952.390 3.670 968.570 4.280 ;
        RECT 969.410 3.670 985.590 4.280 ;
        RECT 986.430 3.670 1002.150 4.280 ;
        RECT 1002.990 3.670 1019.170 4.280 ;
        RECT 1020.010 3.670 1036.190 4.280 ;
        RECT 1037.030 3.670 1052.750 4.280 ;
        RECT 1053.590 3.670 1069.770 4.280 ;
        RECT 1070.610 3.670 1086.330 4.280 ;
        RECT 1087.170 3.670 1103.350 4.280 ;
        RECT 1104.190 3.670 1120.370 4.280 ;
        RECT 1121.210 3.670 1136.930 4.280 ;
        RECT 1137.770 3.670 1153.950 4.280 ;
        RECT 1154.790 3.670 1170.970 4.280 ;
        RECT 1171.810 3.670 1187.530 4.280 ;
        RECT 1188.370 3.670 1204.550 4.280 ;
        RECT 1205.390 3.670 1221.570 4.280 ;
        RECT 1222.410 3.670 1238.130 4.280 ;
        RECT 1238.970 3.670 1255.150 4.280 ;
        RECT 1255.990 3.670 1272.170 4.280 ;
        RECT 1273.010 3.670 1288.730 4.280 ;
        RECT 1289.570 3.670 1305.750 4.280 ;
        RECT 1306.590 3.670 1322.310 4.280 ;
        RECT 1323.150 3.670 1339.330 4.280 ;
        RECT 1340.170 3.670 1356.350 4.280 ;
        RECT 1357.190 3.670 1372.910 4.280 ;
        RECT 1373.750 3.670 1389.930 4.280 ;
        RECT 1390.770 3.670 1406.950 4.280 ;
        RECT 1407.790 3.670 1423.510 4.280 ;
        RECT 1424.350 3.670 1440.530 4.280 ;
        RECT 1441.370 3.670 1457.550 4.280 ;
        RECT 1458.390 3.670 1474.110 4.280 ;
        RECT 1474.950 3.670 1491.130 4.280 ;
        RECT 1491.970 3.670 1493.060 4.280 ;
      LAYER met3 ;
        RECT 4.400 1490.240 1496.000 1490.385 ;
        RECT 4.400 1489.520 1495.600 1490.240 ;
        RECT 4.000 1488.840 1495.600 1489.520 ;
        RECT 4.000 1471.880 1496.000 1488.840 ;
        RECT 4.400 1470.480 1496.000 1471.880 ;
        RECT 4.000 1469.160 1496.000 1470.480 ;
        RECT 4.000 1467.760 1495.600 1469.160 ;
        RECT 4.000 1453.520 1496.000 1467.760 ;
        RECT 4.400 1452.120 1496.000 1453.520 ;
        RECT 4.000 1448.760 1496.000 1452.120 ;
        RECT 4.000 1447.360 1495.600 1448.760 ;
        RECT 4.000 1434.480 1496.000 1447.360 ;
        RECT 4.400 1433.080 1496.000 1434.480 ;
        RECT 4.000 1427.680 1496.000 1433.080 ;
        RECT 4.000 1426.280 1495.600 1427.680 ;
        RECT 4.000 1416.120 1496.000 1426.280 ;
        RECT 4.400 1414.720 1496.000 1416.120 ;
        RECT 4.000 1406.600 1496.000 1414.720 ;
        RECT 4.000 1405.200 1495.600 1406.600 ;
        RECT 4.000 1397.080 1496.000 1405.200 ;
        RECT 4.400 1395.680 1496.000 1397.080 ;
        RECT 4.000 1386.200 1496.000 1395.680 ;
        RECT 4.000 1384.800 1495.600 1386.200 ;
        RECT 4.000 1378.040 1496.000 1384.800 ;
        RECT 4.400 1376.640 1496.000 1378.040 ;
        RECT 4.000 1365.120 1496.000 1376.640 ;
        RECT 4.000 1363.720 1495.600 1365.120 ;
        RECT 4.000 1359.680 1496.000 1363.720 ;
        RECT 4.400 1358.280 1496.000 1359.680 ;
        RECT 4.000 1344.040 1496.000 1358.280 ;
        RECT 4.000 1342.640 1495.600 1344.040 ;
        RECT 4.000 1340.640 1496.000 1342.640 ;
        RECT 4.400 1339.240 1496.000 1340.640 ;
        RECT 4.000 1323.640 1496.000 1339.240 ;
        RECT 4.000 1322.280 1495.600 1323.640 ;
        RECT 4.400 1322.240 1495.600 1322.280 ;
        RECT 4.400 1320.880 1496.000 1322.240 ;
        RECT 4.000 1303.240 1496.000 1320.880 ;
        RECT 4.400 1302.560 1496.000 1303.240 ;
        RECT 4.400 1301.840 1495.600 1302.560 ;
        RECT 4.000 1301.160 1495.600 1301.840 ;
        RECT 4.000 1284.880 1496.000 1301.160 ;
        RECT 4.400 1283.480 1496.000 1284.880 ;
        RECT 4.000 1281.480 1496.000 1283.480 ;
        RECT 4.000 1280.080 1495.600 1281.480 ;
        RECT 4.000 1265.840 1496.000 1280.080 ;
        RECT 4.400 1264.440 1496.000 1265.840 ;
        RECT 4.000 1261.080 1496.000 1264.440 ;
        RECT 4.000 1259.680 1495.600 1261.080 ;
        RECT 4.000 1246.800 1496.000 1259.680 ;
        RECT 4.400 1245.400 1496.000 1246.800 ;
        RECT 4.000 1240.000 1496.000 1245.400 ;
        RECT 4.000 1238.600 1495.600 1240.000 ;
        RECT 4.000 1228.440 1496.000 1238.600 ;
        RECT 4.400 1227.040 1496.000 1228.440 ;
        RECT 4.000 1219.600 1496.000 1227.040 ;
        RECT 4.000 1218.200 1495.600 1219.600 ;
        RECT 4.000 1209.400 1496.000 1218.200 ;
        RECT 4.400 1208.000 1496.000 1209.400 ;
        RECT 4.000 1198.520 1496.000 1208.000 ;
        RECT 4.000 1197.120 1495.600 1198.520 ;
        RECT 4.000 1191.040 1496.000 1197.120 ;
        RECT 4.400 1189.640 1496.000 1191.040 ;
        RECT 4.000 1177.440 1496.000 1189.640 ;
        RECT 4.000 1176.040 1495.600 1177.440 ;
        RECT 4.000 1172.000 1496.000 1176.040 ;
        RECT 4.400 1170.600 1496.000 1172.000 ;
        RECT 4.000 1157.040 1496.000 1170.600 ;
        RECT 4.000 1155.640 1495.600 1157.040 ;
        RECT 4.000 1153.640 1496.000 1155.640 ;
        RECT 4.400 1152.240 1496.000 1153.640 ;
        RECT 4.000 1135.960 1496.000 1152.240 ;
        RECT 4.000 1134.600 1495.600 1135.960 ;
        RECT 4.400 1134.560 1495.600 1134.600 ;
        RECT 4.400 1133.200 1496.000 1134.560 ;
        RECT 4.000 1115.560 1496.000 1133.200 ;
        RECT 4.400 1114.880 1496.000 1115.560 ;
        RECT 4.400 1114.160 1495.600 1114.880 ;
        RECT 4.000 1113.480 1495.600 1114.160 ;
        RECT 4.000 1097.200 1496.000 1113.480 ;
        RECT 4.400 1095.800 1496.000 1097.200 ;
        RECT 4.000 1094.480 1496.000 1095.800 ;
        RECT 4.000 1093.080 1495.600 1094.480 ;
        RECT 4.000 1078.160 1496.000 1093.080 ;
        RECT 4.400 1076.760 1496.000 1078.160 ;
        RECT 4.000 1073.400 1496.000 1076.760 ;
        RECT 4.000 1072.000 1495.600 1073.400 ;
        RECT 4.000 1059.800 1496.000 1072.000 ;
        RECT 4.400 1058.400 1496.000 1059.800 ;
        RECT 4.000 1052.320 1496.000 1058.400 ;
        RECT 4.000 1050.920 1495.600 1052.320 ;
        RECT 4.000 1040.760 1496.000 1050.920 ;
        RECT 4.400 1039.360 1496.000 1040.760 ;
        RECT 4.000 1031.920 1496.000 1039.360 ;
        RECT 4.000 1030.520 1495.600 1031.920 ;
        RECT 4.000 1022.400 1496.000 1030.520 ;
        RECT 4.400 1021.000 1496.000 1022.400 ;
        RECT 4.000 1010.840 1496.000 1021.000 ;
        RECT 4.000 1009.440 1495.600 1010.840 ;
        RECT 4.000 1003.360 1496.000 1009.440 ;
        RECT 4.400 1001.960 1496.000 1003.360 ;
        RECT 4.000 990.440 1496.000 1001.960 ;
        RECT 4.000 989.040 1495.600 990.440 ;
        RECT 4.000 984.320 1496.000 989.040 ;
        RECT 4.400 982.920 1496.000 984.320 ;
        RECT 4.000 969.360 1496.000 982.920 ;
        RECT 4.000 967.960 1495.600 969.360 ;
        RECT 4.000 965.960 1496.000 967.960 ;
        RECT 4.400 964.560 1496.000 965.960 ;
        RECT 4.000 948.280 1496.000 964.560 ;
        RECT 4.000 946.920 1495.600 948.280 ;
        RECT 4.400 946.880 1495.600 946.920 ;
        RECT 4.400 945.520 1496.000 946.880 ;
        RECT 4.000 928.560 1496.000 945.520 ;
        RECT 4.400 927.880 1496.000 928.560 ;
        RECT 4.400 927.160 1495.600 927.880 ;
        RECT 4.000 926.480 1495.600 927.160 ;
        RECT 4.000 909.520 1496.000 926.480 ;
        RECT 4.400 908.120 1496.000 909.520 ;
        RECT 4.000 906.800 1496.000 908.120 ;
        RECT 4.000 905.400 1495.600 906.800 ;
        RECT 4.000 891.160 1496.000 905.400 ;
        RECT 4.400 889.760 1496.000 891.160 ;
        RECT 4.000 885.720 1496.000 889.760 ;
        RECT 4.000 884.320 1495.600 885.720 ;
        RECT 4.000 872.120 1496.000 884.320 ;
        RECT 4.400 870.720 1496.000 872.120 ;
        RECT 4.000 865.320 1496.000 870.720 ;
        RECT 4.000 863.920 1495.600 865.320 ;
        RECT 4.000 853.080 1496.000 863.920 ;
        RECT 4.400 851.680 1496.000 853.080 ;
        RECT 4.000 844.240 1496.000 851.680 ;
        RECT 4.000 842.840 1495.600 844.240 ;
        RECT 4.000 834.720 1496.000 842.840 ;
        RECT 4.400 833.320 1496.000 834.720 ;
        RECT 4.000 823.160 1496.000 833.320 ;
        RECT 4.000 821.760 1495.600 823.160 ;
        RECT 4.000 815.680 1496.000 821.760 ;
        RECT 4.400 814.280 1496.000 815.680 ;
        RECT 4.000 802.760 1496.000 814.280 ;
        RECT 4.000 801.360 1495.600 802.760 ;
        RECT 4.000 797.320 1496.000 801.360 ;
        RECT 4.400 795.920 1496.000 797.320 ;
        RECT 4.000 781.680 1496.000 795.920 ;
        RECT 4.000 780.280 1495.600 781.680 ;
        RECT 4.000 778.280 1496.000 780.280 ;
        RECT 4.400 776.880 1496.000 778.280 ;
        RECT 4.000 761.280 1496.000 776.880 ;
        RECT 4.000 759.920 1495.600 761.280 ;
        RECT 4.400 759.880 1495.600 759.920 ;
        RECT 4.400 758.520 1496.000 759.880 ;
        RECT 4.000 740.880 1496.000 758.520 ;
        RECT 4.400 740.200 1496.000 740.880 ;
        RECT 4.400 739.480 1495.600 740.200 ;
        RECT 4.000 738.800 1495.600 739.480 ;
        RECT 4.000 721.840 1496.000 738.800 ;
        RECT 4.400 720.440 1496.000 721.840 ;
        RECT 4.000 719.120 1496.000 720.440 ;
        RECT 4.000 717.720 1495.600 719.120 ;
        RECT 4.000 703.480 1496.000 717.720 ;
        RECT 4.400 702.080 1496.000 703.480 ;
        RECT 4.000 698.720 1496.000 702.080 ;
        RECT 4.000 697.320 1495.600 698.720 ;
        RECT 4.000 684.440 1496.000 697.320 ;
        RECT 4.400 683.040 1496.000 684.440 ;
        RECT 4.000 677.640 1496.000 683.040 ;
        RECT 4.000 676.240 1495.600 677.640 ;
        RECT 4.000 666.080 1496.000 676.240 ;
        RECT 4.400 664.680 1496.000 666.080 ;
        RECT 4.000 656.560 1496.000 664.680 ;
        RECT 4.000 655.160 1495.600 656.560 ;
        RECT 4.000 647.040 1496.000 655.160 ;
        RECT 4.400 645.640 1496.000 647.040 ;
        RECT 4.000 636.160 1496.000 645.640 ;
        RECT 4.000 634.760 1495.600 636.160 ;
        RECT 4.000 628.000 1496.000 634.760 ;
        RECT 4.400 626.600 1496.000 628.000 ;
        RECT 4.000 615.080 1496.000 626.600 ;
        RECT 4.000 613.680 1495.600 615.080 ;
        RECT 4.000 609.640 1496.000 613.680 ;
        RECT 4.400 608.240 1496.000 609.640 ;
        RECT 4.000 594.000 1496.000 608.240 ;
        RECT 4.000 592.600 1495.600 594.000 ;
        RECT 4.000 590.600 1496.000 592.600 ;
        RECT 4.400 589.200 1496.000 590.600 ;
        RECT 4.000 573.600 1496.000 589.200 ;
        RECT 4.000 572.240 1495.600 573.600 ;
        RECT 4.400 572.200 1495.600 572.240 ;
        RECT 4.400 570.840 1496.000 572.200 ;
        RECT 4.000 553.200 1496.000 570.840 ;
        RECT 4.400 552.520 1496.000 553.200 ;
        RECT 4.400 551.800 1495.600 552.520 ;
        RECT 4.000 551.120 1495.600 551.800 ;
        RECT 4.000 534.840 1496.000 551.120 ;
        RECT 4.400 533.440 1496.000 534.840 ;
        RECT 4.000 531.440 1496.000 533.440 ;
        RECT 4.000 530.040 1495.600 531.440 ;
        RECT 4.000 515.800 1496.000 530.040 ;
        RECT 4.400 514.400 1496.000 515.800 ;
        RECT 4.000 511.040 1496.000 514.400 ;
        RECT 4.000 509.640 1495.600 511.040 ;
        RECT 4.000 496.760 1496.000 509.640 ;
        RECT 4.400 495.360 1496.000 496.760 ;
        RECT 4.000 489.960 1496.000 495.360 ;
        RECT 4.000 488.560 1495.600 489.960 ;
        RECT 4.000 478.400 1496.000 488.560 ;
        RECT 4.400 477.000 1496.000 478.400 ;
        RECT 4.000 469.560 1496.000 477.000 ;
        RECT 4.000 468.160 1495.600 469.560 ;
        RECT 4.000 459.360 1496.000 468.160 ;
        RECT 4.400 457.960 1496.000 459.360 ;
        RECT 4.000 448.480 1496.000 457.960 ;
        RECT 4.000 447.080 1495.600 448.480 ;
        RECT 4.000 441.000 1496.000 447.080 ;
        RECT 4.400 439.600 1496.000 441.000 ;
        RECT 4.000 427.400 1496.000 439.600 ;
        RECT 4.000 426.000 1495.600 427.400 ;
        RECT 4.000 421.960 1496.000 426.000 ;
        RECT 4.400 420.560 1496.000 421.960 ;
        RECT 4.000 407.000 1496.000 420.560 ;
        RECT 4.000 405.600 1495.600 407.000 ;
        RECT 4.000 403.600 1496.000 405.600 ;
        RECT 4.400 402.200 1496.000 403.600 ;
        RECT 4.000 385.920 1496.000 402.200 ;
        RECT 4.000 384.560 1495.600 385.920 ;
        RECT 4.400 384.520 1495.600 384.560 ;
        RECT 4.400 383.160 1496.000 384.520 ;
        RECT 4.000 365.520 1496.000 383.160 ;
        RECT 4.400 364.840 1496.000 365.520 ;
        RECT 4.400 364.120 1495.600 364.840 ;
        RECT 4.000 363.440 1495.600 364.120 ;
        RECT 4.000 347.160 1496.000 363.440 ;
        RECT 4.400 345.760 1496.000 347.160 ;
        RECT 4.000 344.440 1496.000 345.760 ;
        RECT 4.000 343.040 1495.600 344.440 ;
        RECT 4.000 328.120 1496.000 343.040 ;
        RECT 4.400 326.720 1496.000 328.120 ;
        RECT 4.000 323.360 1496.000 326.720 ;
        RECT 4.000 321.960 1495.600 323.360 ;
        RECT 4.000 309.760 1496.000 321.960 ;
        RECT 4.400 308.360 1496.000 309.760 ;
        RECT 4.000 302.280 1496.000 308.360 ;
        RECT 4.000 300.880 1495.600 302.280 ;
        RECT 4.000 290.720 1496.000 300.880 ;
        RECT 4.400 289.320 1496.000 290.720 ;
        RECT 4.000 281.880 1496.000 289.320 ;
        RECT 4.000 280.480 1495.600 281.880 ;
        RECT 4.000 272.360 1496.000 280.480 ;
        RECT 4.400 270.960 1496.000 272.360 ;
        RECT 4.000 260.800 1496.000 270.960 ;
        RECT 4.000 259.400 1495.600 260.800 ;
        RECT 4.000 253.320 1496.000 259.400 ;
        RECT 4.400 251.920 1496.000 253.320 ;
        RECT 4.000 240.400 1496.000 251.920 ;
        RECT 4.000 239.000 1495.600 240.400 ;
        RECT 4.000 234.280 1496.000 239.000 ;
        RECT 4.400 232.880 1496.000 234.280 ;
        RECT 4.000 219.320 1496.000 232.880 ;
        RECT 4.000 217.920 1495.600 219.320 ;
        RECT 4.000 215.920 1496.000 217.920 ;
        RECT 4.400 214.520 1496.000 215.920 ;
        RECT 4.000 198.240 1496.000 214.520 ;
        RECT 4.000 196.880 1495.600 198.240 ;
        RECT 4.400 196.840 1495.600 196.880 ;
        RECT 4.400 195.480 1496.000 196.840 ;
        RECT 4.000 178.520 1496.000 195.480 ;
        RECT 4.400 177.840 1496.000 178.520 ;
        RECT 4.400 177.120 1495.600 177.840 ;
        RECT 4.000 176.440 1495.600 177.120 ;
        RECT 4.000 159.480 1496.000 176.440 ;
        RECT 4.400 158.080 1496.000 159.480 ;
        RECT 4.000 156.760 1496.000 158.080 ;
        RECT 4.000 155.360 1495.600 156.760 ;
        RECT 4.000 141.120 1496.000 155.360 ;
        RECT 4.400 139.720 1496.000 141.120 ;
        RECT 4.000 135.680 1496.000 139.720 ;
        RECT 4.000 134.280 1495.600 135.680 ;
        RECT 4.000 122.080 1496.000 134.280 ;
        RECT 4.400 120.680 1496.000 122.080 ;
        RECT 4.000 115.280 1496.000 120.680 ;
        RECT 4.000 113.880 1495.600 115.280 ;
        RECT 4.000 103.040 1496.000 113.880 ;
        RECT 4.400 101.640 1496.000 103.040 ;
        RECT 4.000 94.200 1496.000 101.640 ;
        RECT 4.000 92.800 1495.600 94.200 ;
        RECT 4.000 84.680 1496.000 92.800 ;
        RECT 4.400 83.280 1496.000 84.680 ;
        RECT 4.000 73.120 1496.000 83.280 ;
        RECT 4.000 71.720 1495.600 73.120 ;
        RECT 4.000 65.640 1496.000 71.720 ;
        RECT 4.400 64.240 1496.000 65.640 ;
        RECT 4.000 52.720 1496.000 64.240 ;
        RECT 4.000 51.320 1495.600 52.720 ;
        RECT 4.000 47.280 1496.000 51.320 ;
        RECT 4.400 45.880 1496.000 47.280 ;
        RECT 4.000 31.640 1496.000 45.880 ;
        RECT 4.000 30.240 1495.600 31.640 ;
        RECT 4.000 28.240 1496.000 30.240 ;
        RECT 4.400 26.840 1496.000 28.240 ;
        RECT 4.000 11.240 1496.000 26.840 ;
        RECT 4.000 9.880 1495.600 11.240 ;
        RECT 4.400 9.840 1495.600 9.880 ;
        RECT 4.400 9.015 1496.000 9.840 ;
      LAYER met4 ;
        RECT 96.895 11.735 97.440 1485.625 ;
        RECT 99.840 11.735 174.240 1485.625 ;
        RECT 176.640 11.735 251.040 1485.625 ;
        RECT 253.440 11.735 327.840 1485.625 ;
        RECT 330.240 11.735 404.640 1485.625 ;
        RECT 407.040 11.735 481.440 1485.625 ;
        RECT 483.840 11.735 558.240 1485.625 ;
        RECT 560.640 11.735 635.040 1485.625 ;
        RECT 637.440 11.735 711.840 1485.625 ;
        RECT 714.240 11.735 788.640 1485.625 ;
        RECT 791.040 11.735 865.440 1485.625 ;
        RECT 867.840 11.735 942.240 1485.625 ;
        RECT 944.640 11.735 962.945 1485.625 ;
  END
END core
END LIBRARY

