VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 1496.000 104.790 1500.000 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1311.760 1500.000 1312.360 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.130 0.000 1184.410 4.000 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.630 0.000 1218.910 4.000 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1334.200 4.000 1334.800 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 1496.000 1298.490 1500.000 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 0.000 1269.970 4.000 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.730 0.000 1304.010 4.000 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 0.000 1321.030 4.000 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 1496.000 346.750 1500.000 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1372.960 4.000 1373.560 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1360.720 1500.000 1361.320 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.770 0.000 1338.050 4.000 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.720 4.000 1412.320 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1377.040 1500.000 1377.640 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 0.000 1406.130 4.000 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.610 1496.000 1362.890 1500.000 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.910 0.000 1457.190 4.000 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.160 4.000 1451.760 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.920 4.000 1490.520 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1393.360 1500.000 1393.960 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 1496.000 1427.290 1500.000 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 0.000 1474.210 4.000 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.210 1496.000 1459.490 1500.000 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 1496.000 1475.590 1500.000 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 1496.000 1491.690 1500.000 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1474.960 1500.000 1475.560 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 235.320 1500.000 235.920 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 300.600 1500.000 301.200 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 333.240 1500.000 333.840 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 398.520 1500.000 399.120 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 463.800 1500.000 464.400 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 1496.000 153.090 1500.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 496.440 1500.000 497.040 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 561.720 1500.000 562.320 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 1496.000 572.610 1500.000 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 1496.000 620.910 1500.000 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 692.280 1500.000 692.880 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 1496.000 201.390 1500.000 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 741.240 1500.000 741.840 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 1496.000 669.210 1500.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 789.520 1500.000 790.120 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 805.840 1500.000 806.440 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 822.160 1500.000 822.760 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 854.800 1500.000 855.400 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 871.120 1500.000 871.720 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 55.800 1500.000 56.400 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 1496.000 733.610 1500.000 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 0.000 639.310 4.000 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.160 4.000 788.760 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 1496.000 782.370 1500.000 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 4.000 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 1496.000 814.570 1500.000 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 4.000 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 0.000 809.510 4.000 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 920.080 1500.000 920.680 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 1496.000 878.970 1500.000 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.120 4.000 905.720 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 1496.000 911.170 1500.000 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 952.720 1500.000 953.320 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 969.040 1500.000 969.640 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 1496.000 943.370 1500.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 0.000 912.090 4.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.800 4.000 1042.400 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1061.520 4.000 1062.120 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1080.560 4.000 1081.160 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 1496.000 282.350 1500.000 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.850 0.000 946.130 4.000 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1100.280 4.000 1100.880 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1066.960 1500.000 1067.560 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1099.600 1500.000 1100.200 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1115.920 1500.000 1116.520 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 1496.000 975.570 1500.000 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 1496.000 991.670 1500.000 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1158.760 4.000 1159.360 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 0.000 1014.210 4.000 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1496.000 1008.230 1500.000 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1164.880 1500.000 1165.480 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1496.000 1040.430 1500.000 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 1496.000 1056.530 1500.000 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 0.000 1048.250 4.000 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.280 4.000 1236.880 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 0.000 1065.270 4.000 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1197.520 1500.000 1198.120 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1213.840 1500.000 1214.440 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 1496.000 1104.830 1500.000 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 1496.000 1120.930 1500.000 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 1496.000 1137.030 1500.000 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.720 4.000 1276.320 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 1496.000 1153.130 1500.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1294.760 4.000 1295.360 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 1496.000 1185.330 1500.000 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1314.480 4.000 1315.080 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.110 0.000 1167.390 4.000 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1279.120 1500.000 1279.720 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1496.000 1217.530 1500.000 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 251.640 1500.000 252.240 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 1496.000 378.950 1500.000 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 349.560 1500.000 350.160 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 414.840 1500.000 415.440 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 447.480 1500.000 448.080 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 1496.000 491.650 1500.000 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 23.160 1500.000 23.760 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 512.760 1500.000 513.360 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 610.680 1500.000 611.280 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 1496.000 637.010 1500.000 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 675.960 1500.000 676.560 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 708.600 1500.000 709.200 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 757.560 1500.000 758.160 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 1496.000 233.590 1500.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 1496.000 298.450 1500.000 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 202.680 1500.000 203.280 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 1496.000 40.390 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 1496.000 88.690 1500.000 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 1496.000 72.590 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 1496.000 56.490 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 7.520 1500.000 8.120 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 219.000 1500.000 219.600 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 267.960 1500.000 268.560 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 316.920 1500.000 317.520 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 365.880 1500.000 366.480 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 1496.000 427.250 1500.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 431.160 1500.000 431.760 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 1496.000 169.190 1500.000 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 72.120 1500.000 72.720 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 1496.000 249.690 1500.000 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 121.080 1500.000 121.680 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 1496.000 330.650 1500.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 1496.000 120.890 1500.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 1496.000 1249.730 1500.000 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 1496.000 1266.290 1500.000 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.110 1496.000 1282.390 1500.000 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.650 0.000 1235.930 4.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 1496.000 1314.590 1500.000 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.710 0.000 1286.990 4.000 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1328.080 1500.000 1328.680 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 1496.000 1330.690 1500.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1344.400 1500.000 1345.000 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.510 1496.000 1346.790 1500.000 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.680 4.000 1393.280 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.790 0.000 1355.070 4.000 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 0.000 1372.090 4.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.830 0.000 1389.110 4.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 0.000 1440.170 4.000 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 1496.000 1378.990 1500.000 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.810 1496.000 1395.090 1500.000 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1470.200 4.000 1470.800 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 1496.000 1411.190 1500.000 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1409.680 1500.000 1410.280 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.110 1496.000 1443.390 1500.000 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1426.000 1500.000 1426.600 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1442.320 1500.000 1442.920 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1458.640 1500.000 1459.240 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1491.280 1500.000 1491.880 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 284.280 1500.000 284.880 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 1496.000 395.050 1500.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 382.200 1500.000 382.800 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 1496.000 459.450 1500.000 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 1496.000 524.310 1500.000 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 1496.000 185.290 1500.000 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 480.120 1500.000 480.720 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 1496.000 556.510 1500.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 529.080 1500.000 529.680 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 578.040 1500.000 578.640 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 1496.000 588.710 1500.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 4.000 594.280 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 643.320 1500.000 643.920 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 659.640 1500.000 660.240 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 1496.000 653.110 1500.000 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 1496.000 217.490 1500.000 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 773.200 1500.000 773.800 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 1496.000 685.310 1500.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 1496.000 701.410 1500.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 838.480 1500.000 839.080 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 1496.000 717.510 1500.000 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 88.440 1500.000 89.040 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.120 4.000 769.720 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 1496.000 749.710 1500.000 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 887.440 1500.000 888.040 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 1496.000 766.270 1500.000 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 903.760 1500.000 904.360 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 1496.000 798.470 1500.000 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 827.600 4.000 828.200 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 1496.000 830.670 1500.000 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 1496.000 846.770 1500.000 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 1496.000 862.870 1500.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 4.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 0.000 877.590 4.000 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 936.400 1500.000 937.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 1496.000 895.070 1500.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 137.400 1500.000 138.000 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 944.560 4.000 945.160 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 963.600 4.000 964.200 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 0.000 894.610 4.000 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 1496.000 927.270 1500.000 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 985.360 1500.000 985.960 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1022.080 4.000 1022.680 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 1496.000 959.470 1500.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1001.680 1500.000 1002.280 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1018.000 1500.000 1018.600 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 0.000 929.110 4.000 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 1496.000 314.550 1500.000 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1034.320 1500.000 1034.920 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1050.640 1500.000 1051.240 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1083.280 1500.000 1083.880 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.000 4.000 1120.600 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1132.240 1500.000 1132.840 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 0.000 980.170 4.000 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 0.000 997.190 4.000 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.800 4.000 1178.400 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1148.560 1500.000 1149.160 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 153.720 1500.000 154.320 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1197.520 4.000 1198.120 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 1496.000 1024.330 1500.000 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 0.000 1031.230 4.000 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1181.200 1500.000 1181.800 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.240 4.000 1217.840 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1496.000 1072.630 1500.000 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 1496.000 1088.730 1500.000 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 0.000 1099.310 4.000 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1230.160 1500.000 1230.760 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 186.360 1500.000 186.960 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.050 0.000 1116.330 4.000 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1256.000 4.000 1256.600 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.070 0.000 1133.350 4.000 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 1496.000 1169.230 1500.000 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1246.480 1500.000 1247.080 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 0.000 1150.370 4.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1262.800 1500.000 1263.400 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 1496.000 1201.430 1500.000 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1295.440 1500.000 1296.040 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1496.000 1233.630 1500.000 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 1496.000 8.190 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 1496.000 24.290 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 1496.000 136.990 1500.000 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 1496.000 362.850 1500.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 1496.000 411.150 1500.000 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 1496.000 443.350 1500.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 1496.000 475.550 1500.000 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 1496.000 508.210 1500.000 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 1496.000 540.410 1500.000 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 545.400 1500.000 546.000 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 594.360 1500.000 594.960 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1496.000 604.810 1500.000 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 627.000 1500.000 627.600 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 724.920 1500.000 725.520 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 39.480 1500.000 40.080 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 104.760 1500.000 105.360 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 1496.000 266.250 1500.000 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 170.040 1500.000 170.640 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.080 1488.080 ;
      LAYER met2 ;
        RECT 6.990 1495.720 7.630 1496.410 ;
        RECT 8.470 1495.720 23.730 1496.410 ;
        RECT 24.570 1495.720 39.830 1496.410 ;
        RECT 40.670 1495.720 55.930 1496.410 ;
        RECT 56.770 1495.720 72.030 1496.410 ;
        RECT 72.870 1495.720 88.130 1496.410 ;
        RECT 88.970 1495.720 104.230 1496.410 ;
        RECT 105.070 1495.720 120.330 1496.410 ;
        RECT 121.170 1495.720 136.430 1496.410 ;
        RECT 137.270 1495.720 152.530 1496.410 ;
        RECT 153.370 1495.720 168.630 1496.410 ;
        RECT 169.470 1495.720 184.730 1496.410 ;
        RECT 185.570 1495.720 200.830 1496.410 ;
        RECT 201.670 1495.720 216.930 1496.410 ;
        RECT 217.770 1495.720 233.030 1496.410 ;
        RECT 233.870 1495.720 249.130 1496.410 ;
        RECT 249.970 1495.720 265.690 1496.410 ;
        RECT 266.530 1495.720 281.790 1496.410 ;
        RECT 282.630 1495.720 297.890 1496.410 ;
        RECT 298.730 1495.720 313.990 1496.410 ;
        RECT 314.830 1495.720 330.090 1496.410 ;
        RECT 330.930 1495.720 346.190 1496.410 ;
        RECT 347.030 1495.720 362.290 1496.410 ;
        RECT 363.130 1495.720 378.390 1496.410 ;
        RECT 379.230 1495.720 394.490 1496.410 ;
        RECT 395.330 1495.720 410.590 1496.410 ;
        RECT 411.430 1495.720 426.690 1496.410 ;
        RECT 427.530 1495.720 442.790 1496.410 ;
        RECT 443.630 1495.720 458.890 1496.410 ;
        RECT 459.730 1495.720 474.990 1496.410 ;
        RECT 475.830 1495.720 491.090 1496.410 ;
        RECT 491.930 1495.720 507.650 1496.410 ;
        RECT 508.490 1495.720 523.750 1496.410 ;
        RECT 524.590 1495.720 539.850 1496.410 ;
        RECT 540.690 1495.720 555.950 1496.410 ;
        RECT 556.790 1495.720 572.050 1496.410 ;
        RECT 572.890 1495.720 588.150 1496.410 ;
        RECT 588.990 1495.720 604.250 1496.410 ;
        RECT 605.090 1495.720 620.350 1496.410 ;
        RECT 621.190 1495.720 636.450 1496.410 ;
        RECT 637.290 1495.720 652.550 1496.410 ;
        RECT 653.390 1495.720 668.650 1496.410 ;
        RECT 669.490 1495.720 684.750 1496.410 ;
        RECT 685.590 1495.720 700.850 1496.410 ;
        RECT 701.690 1495.720 716.950 1496.410 ;
        RECT 717.790 1495.720 733.050 1496.410 ;
        RECT 733.890 1495.720 749.150 1496.410 ;
        RECT 749.990 1495.720 765.710 1496.410 ;
        RECT 766.550 1495.720 781.810 1496.410 ;
        RECT 782.650 1495.720 797.910 1496.410 ;
        RECT 798.750 1495.720 814.010 1496.410 ;
        RECT 814.850 1495.720 830.110 1496.410 ;
        RECT 830.950 1495.720 846.210 1496.410 ;
        RECT 847.050 1495.720 862.310 1496.410 ;
        RECT 863.150 1495.720 878.410 1496.410 ;
        RECT 879.250 1495.720 894.510 1496.410 ;
        RECT 895.350 1495.720 910.610 1496.410 ;
        RECT 911.450 1495.720 926.710 1496.410 ;
        RECT 927.550 1495.720 942.810 1496.410 ;
        RECT 943.650 1495.720 958.910 1496.410 ;
        RECT 959.750 1495.720 975.010 1496.410 ;
        RECT 975.850 1495.720 991.110 1496.410 ;
        RECT 991.950 1495.720 1007.670 1496.410 ;
        RECT 1008.510 1495.720 1023.770 1496.410 ;
        RECT 1024.610 1495.720 1039.870 1496.410 ;
        RECT 1040.710 1495.720 1055.970 1496.410 ;
        RECT 1056.810 1495.720 1072.070 1496.410 ;
        RECT 1072.910 1495.720 1088.170 1496.410 ;
        RECT 1089.010 1495.720 1104.270 1496.410 ;
        RECT 1105.110 1495.720 1120.370 1496.410 ;
        RECT 1121.210 1495.720 1136.470 1496.410 ;
        RECT 1137.310 1495.720 1152.570 1496.410 ;
        RECT 1153.410 1495.720 1168.670 1496.410 ;
        RECT 1169.510 1495.720 1184.770 1496.410 ;
        RECT 1185.610 1495.720 1200.870 1496.410 ;
        RECT 1201.710 1495.720 1216.970 1496.410 ;
        RECT 1217.810 1495.720 1233.070 1496.410 ;
        RECT 1233.910 1495.720 1249.170 1496.410 ;
        RECT 1250.010 1495.720 1265.730 1496.410 ;
        RECT 1266.570 1495.720 1281.830 1496.410 ;
        RECT 1282.670 1495.720 1297.930 1496.410 ;
        RECT 1298.770 1495.720 1314.030 1496.410 ;
        RECT 1314.870 1495.720 1330.130 1496.410 ;
        RECT 1330.970 1495.720 1346.230 1496.410 ;
        RECT 1347.070 1495.720 1362.330 1496.410 ;
        RECT 1363.170 1495.720 1378.430 1496.410 ;
        RECT 1379.270 1495.720 1394.530 1496.410 ;
        RECT 1395.370 1495.720 1410.630 1496.410 ;
        RECT 1411.470 1495.720 1426.730 1496.410 ;
        RECT 1427.570 1495.720 1442.830 1496.410 ;
        RECT 1443.670 1495.720 1458.930 1496.410 ;
        RECT 1459.770 1495.720 1475.030 1496.410 ;
        RECT 1475.870 1495.720 1491.130 1496.410 ;
        RECT 6.990 4.280 1491.680 1495.720 ;
        RECT 6.990 3.670 8.090 4.280 ;
        RECT 8.930 3.670 25.110 4.280 ;
        RECT 25.950 3.670 42.130 4.280 ;
        RECT 42.970 3.670 59.150 4.280 ;
        RECT 59.990 3.670 76.170 4.280 ;
        RECT 77.010 3.670 93.190 4.280 ;
        RECT 94.030 3.670 110.210 4.280 ;
        RECT 111.050 3.670 127.230 4.280 ;
        RECT 128.070 3.670 144.250 4.280 ;
        RECT 145.090 3.670 161.270 4.280 ;
        RECT 162.110 3.670 178.290 4.280 ;
        RECT 179.130 3.670 195.310 4.280 ;
        RECT 196.150 3.670 212.330 4.280 ;
        RECT 213.170 3.670 229.350 4.280 ;
        RECT 230.190 3.670 246.370 4.280 ;
        RECT 247.210 3.670 263.390 4.280 ;
        RECT 264.230 3.670 280.410 4.280 ;
        RECT 281.250 3.670 297.430 4.280 ;
        RECT 298.270 3.670 314.910 4.280 ;
        RECT 315.750 3.670 331.930 4.280 ;
        RECT 332.770 3.670 348.950 4.280 ;
        RECT 349.790 3.670 365.970 4.280 ;
        RECT 366.810 3.670 382.990 4.280 ;
        RECT 383.830 3.670 400.010 4.280 ;
        RECT 400.850 3.670 417.030 4.280 ;
        RECT 417.870 3.670 434.050 4.280 ;
        RECT 434.890 3.670 451.070 4.280 ;
        RECT 451.910 3.670 468.090 4.280 ;
        RECT 468.930 3.670 485.110 4.280 ;
        RECT 485.950 3.670 502.130 4.280 ;
        RECT 502.970 3.670 519.150 4.280 ;
        RECT 519.990 3.670 536.170 4.280 ;
        RECT 537.010 3.670 553.190 4.280 ;
        RECT 554.030 3.670 570.210 4.280 ;
        RECT 571.050 3.670 587.230 4.280 ;
        RECT 588.070 3.670 604.250 4.280 ;
        RECT 605.090 3.670 621.730 4.280 ;
        RECT 622.570 3.670 638.750 4.280 ;
        RECT 639.590 3.670 655.770 4.280 ;
        RECT 656.610 3.670 672.790 4.280 ;
        RECT 673.630 3.670 689.810 4.280 ;
        RECT 690.650 3.670 706.830 4.280 ;
        RECT 707.670 3.670 723.850 4.280 ;
        RECT 724.690 3.670 740.870 4.280 ;
        RECT 741.710 3.670 757.890 4.280 ;
        RECT 758.730 3.670 774.910 4.280 ;
        RECT 775.750 3.670 791.930 4.280 ;
        RECT 792.770 3.670 808.950 4.280 ;
        RECT 809.790 3.670 825.970 4.280 ;
        RECT 826.810 3.670 842.990 4.280 ;
        RECT 843.830 3.670 860.010 4.280 ;
        RECT 860.850 3.670 877.030 4.280 ;
        RECT 877.870 3.670 894.050 4.280 ;
        RECT 894.890 3.670 911.530 4.280 ;
        RECT 912.370 3.670 928.550 4.280 ;
        RECT 929.390 3.670 945.570 4.280 ;
        RECT 946.410 3.670 962.590 4.280 ;
        RECT 963.430 3.670 979.610 4.280 ;
        RECT 980.450 3.670 996.630 4.280 ;
        RECT 997.470 3.670 1013.650 4.280 ;
        RECT 1014.490 3.670 1030.670 4.280 ;
        RECT 1031.510 3.670 1047.690 4.280 ;
        RECT 1048.530 3.670 1064.710 4.280 ;
        RECT 1065.550 3.670 1081.730 4.280 ;
        RECT 1082.570 3.670 1098.750 4.280 ;
        RECT 1099.590 3.670 1115.770 4.280 ;
        RECT 1116.610 3.670 1132.790 4.280 ;
        RECT 1133.630 3.670 1149.810 4.280 ;
        RECT 1150.650 3.670 1166.830 4.280 ;
        RECT 1167.670 3.670 1183.850 4.280 ;
        RECT 1184.690 3.670 1200.870 4.280 ;
        RECT 1201.710 3.670 1218.350 4.280 ;
        RECT 1219.190 3.670 1235.370 4.280 ;
        RECT 1236.210 3.670 1252.390 4.280 ;
        RECT 1253.230 3.670 1269.410 4.280 ;
        RECT 1270.250 3.670 1286.430 4.280 ;
        RECT 1287.270 3.670 1303.450 4.280 ;
        RECT 1304.290 3.670 1320.470 4.280 ;
        RECT 1321.310 3.670 1337.490 4.280 ;
        RECT 1338.330 3.670 1354.510 4.280 ;
        RECT 1355.350 3.670 1371.530 4.280 ;
        RECT 1372.370 3.670 1388.550 4.280 ;
        RECT 1389.390 3.670 1405.570 4.280 ;
        RECT 1406.410 3.670 1422.590 4.280 ;
        RECT 1423.430 3.670 1439.610 4.280 ;
        RECT 1440.450 3.670 1456.630 4.280 ;
        RECT 1457.470 3.670 1473.650 4.280 ;
        RECT 1474.490 3.670 1490.670 4.280 ;
        RECT 1491.510 3.670 1491.680 4.280 ;
      LAYER met3 ;
        RECT 4.000 1490.920 1495.600 1491.745 ;
        RECT 4.400 1490.880 1495.600 1490.920 ;
        RECT 4.400 1489.520 1496.000 1490.880 ;
        RECT 4.000 1475.960 1496.000 1489.520 ;
        RECT 4.000 1474.560 1495.600 1475.960 ;
        RECT 4.000 1471.200 1496.000 1474.560 ;
        RECT 4.400 1469.800 1496.000 1471.200 ;
        RECT 4.000 1459.640 1496.000 1469.800 ;
        RECT 4.000 1458.240 1495.600 1459.640 ;
        RECT 4.000 1452.160 1496.000 1458.240 ;
        RECT 4.400 1450.760 1496.000 1452.160 ;
        RECT 4.000 1443.320 1496.000 1450.760 ;
        RECT 4.000 1441.920 1495.600 1443.320 ;
        RECT 4.000 1432.440 1496.000 1441.920 ;
        RECT 4.400 1431.040 1496.000 1432.440 ;
        RECT 4.000 1427.000 1496.000 1431.040 ;
        RECT 4.000 1425.600 1495.600 1427.000 ;
        RECT 4.000 1412.720 1496.000 1425.600 ;
        RECT 4.400 1411.320 1496.000 1412.720 ;
        RECT 4.000 1410.680 1496.000 1411.320 ;
        RECT 4.000 1409.280 1495.600 1410.680 ;
        RECT 4.000 1394.360 1496.000 1409.280 ;
        RECT 4.000 1393.680 1495.600 1394.360 ;
        RECT 4.400 1392.960 1495.600 1393.680 ;
        RECT 4.400 1392.280 1496.000 1392.960 ;
        RECT 4.000 1378.040 1496.000 1392.280 ;
        RECT 4.000 1376.640 1495.600 1378.040 ;
        RECT 4.000 1373.960 1496.000 1376.640 ;
        RECT 4.400 1372.560 1496.000 1373.960 ;
        RECT 4.000 1361.720 1496.000 1372.560 ;
        RECT 4.000 1360.320 1495.600 1361.720 ;
        RECT 4.000 1354.240 1496.000 1360.320 ;
        RECT 4.400 1352.840 1496.000 1354.240 ;
        RECT 4.000 1345.400 1496.000 1352.840 ;
        RECT 4.000 1344.000 1495.600 1345.400 ;
        RECT 4.000 1335.200 1496.000 1344.000 ;
        RECT 4.400 1333.800 1496.000 1335.200 ;
        RECT 4.000 1329.080 1496.000 1333.800 ;
        RECT 4.000 1327.680 1495.600 1329.080 ;
        RECT 4.000 1315.480 1496.000 1327.680 ;
        RECT 4.400 1314.080 1496.000 1315.480 ;
        RECT 4.000 1312.760 1496.000 1314.080 ;
        RECT 4.000 1311.360 1495.600 1312.760 ;
        RECT 4.000 1296.440 1496.000 1311.360 ;
        RECT 4.000 1295.760 1495.600 1296.440 ;
        RECT 4.400 1295.040 1495.600 1295.760 ;
        RECT 4.400 1294.360 1496.000 1295.040 ;
        RECT 4.000 1280.120 1496.000 1294.360 ;
        RECT 4.000 1278.720 1495.600 1280.120 ;
        RECT 4.000 1276.720 1496.000 1278.720 ;
        RECT 4.400 1275.320 1496.000 1276.720 ;
        RECT 4.000 1263.800 1496.000 1275.320 ;
        RECT 4.000 1262.400 1495.600 1263.800 ;
        RECT 4.000 1257.000 1496.000 1262.400 ;
        RECT 4.400 1255.600 1496.000 1257.000 ;
        RECT 4.000 1247.480 1496.000 1255.600 ;
        RECT 4.000 1246.080 1495.600 1247.480 ;
        RECT 4.000 1237.280 1496.000 1246.080 ;
        RECT 4.400 1235.880 1496.000 1237.280 ;
        RECT 4.000 1231.160 1496.000 1235.880 ;
        RECT 4.000 1229.760 1495.600 1231.160 ;
        RECT 4.000 1218.240 1496.000 1229.760 ;
        RECT 4.400 1216.840 1496.000 1218.240 ;
        RECT 4.000 1214.840 1496.000 1216.840 ;
        RECT 4.000 1213.440 1495.600 1214.840 ;
        RECT 4.000 1198.520 1496.000 1213.440 ;
        RECT 4.400 1197.120 1495.600 1198.520 ;
        RECT 4.000 1182.200 1496.000 1197.120 ;
        RECT 4.000 1180.800 1495.600 1182.200 ;
        RECT 4.000 1178.800 1496.000 1180.800 ;
        RECT 4.400 1177.400 1496.000 1178.800 ;
        RECT 4.000 1165.880 1496.000 1177.400 ;
        RECT 4.000 1164.480 1495.600 1165.880 ;
        RECT 4.000 1159.760 1496.000 1164.480 ;
        RECT 4.400 1158.360 1496.000 1159.760 ;
        RECT 4.000 1149.560 1496.000 1158.360 ;
        RECT 4.000 1148.160 1495.600 1149.560 ;
        RECT 4.000 1140.040 1496.000 1148.160 ;
        RECT 4.400 1138.640 1496.000 1140.040 ;
        RECT 4.000 1133.240 1496.000 1138.640 ;
        RECT 4.000 1131.840 1495.600 1133.240 ;
        RECT 4.000 1121.000 1496.000 1131.840 ;
        RECT 4.400 1119.600 1496.000 1121.000 ;
        RECT 4.000 1116.920 1496.000 1119.600 ;
        RECT 4.000 1115.520 1495.600 1116.920 ;
        RECT 4.000 1101.280 1496.000 1115.520 ;
        RECT 4.400 1100.600 1496.000 1101.280 ;
        RECT 4.400 1099.880 1495.600 1100.600 ;
        RECT 4.000 1099.200 1495.600 1099.880 ;
        RECT 4.000 1084.280 1496.000 1099.200 ;
        RECT 4.000 1082.880 1495.600 1084.280 ;
        RECT 4.000 1081.560 1496.000 1082.880 ;
        RECT 4.400 1080.160 1496.000 1081.560 ;
        RECT 4.000 1067.960 1496.000 1080.160 ;
        RECT 4.000 1066.560 1495.600 1067.960 ;
        RECT 4.000 1062.520 1496.000 1066.560 ;
        RECT 4.400 1061.120 1496.000 1062.520 ;
        RECT 4.000 1051.640 1496.000 1061.120 ;
        RECT 4.000 1050.240 1495.600 1051.640 ;
        RECT 4.000 1042.800 1496.000 1050.240 ;
        RECT 4.400 1041.400 1496.000 1042.800 ;
        RECT 4.000 1035.320 1496.000 1041.400 ;
        RECT 4.000 1033.920 1495.600 1035.320 ;
        RECT 4.000 1023.080 1496.000 1033.920 ;
        RECT 4.400 1021.680 1496.000 1023.080 ;
        RECT 4.000 1019.000 1496.000 1021.680 ;
        RECT 4.000 1017.600 1495.600 1019.000 ;
        RECT 4.000 1004.040 1496.000 1017.600 ;
        RECT 4.400 1002.680 1496.000 1004.040 ;
        RECT 4.400 1002.640 1495.600 1002.680 ;
        RECT 4.000 1001.280 1495.600 1002.640 ;
        RECT 4.000 986.360 1496.000 1001.280 ;
        RECT 4.000 984.960 1495.600 986.360 ;
        RECT 4.000 984.320 1496.000 984.960 ;
        RECT 4.400 982.920 1496.000 984.320 ;
        RECT 4.000 970.040 1496.000 982.920 ;
        RECT 4.000 968.640 1495.600 970.040 ;
        RECT 4.000 964.600 1496.000 968.640 ;
        RECT 4.400 963.200 1496.000 964.600 ;
        RECT 4.000 953.720 1496.000 963.200 ;
        RECT 4.000 952.320 1495.600 953.720 ;
        RECT 4.000 945.560 1496.000 952.320 ;
        RECT 4.400 944.160 1496.000 945.560 ;
        RECT 4.000 937.400 1496.000 944.160 ;
        RECT 4.000 936.000 1495.600 937.400 ;
        RECT 4.000 925.840 1496.000 936.000 ;
        RECT 4.400 924.440 1496.000 925.840 ;
        RECT 4.000 921.080 1496.000 924.440 ;
        RECT 4.000 919.680 1495.600 921.080 ;
        RECT 4.000 906.120 1496.000 919.680 ;
        RECT 4.400 904.760 1496.000 906.120 ;
        RECT 4.400 904.720 1495.600 904.760 ;
        RECT 4.000 903.360 1495.600 904.720 ;
        RECT 4.000 888.440 1496.000 903.360 ;
        RECT 4.000 887.080 1495.600 888.440 ;
        RECT 4.400 887.040 1495.600 887.080 ;
        RECT 4.400 885.680 1496.000 887.040 ;
        RECT 4.000 872.120 1496.000 885.680 ;
        RECT 4.000 870.720 1495.600 872.120 ;
        RECT 4.000 867.360 1496.000 870.720 ;
        RECT 4.400 865.960 1496.000 867.360 ;
        RECT 4.000 855.800 1496.000 865.960 ;
        RECT 4.000 854.400 1495.600 855.800 ;
        RECT 4.000 847.640 1496.000 854.400 ;
        RECT 4.400 846.240 1496.000 847.640 ;
        RECT 4.000 839.480 1496.000 846.240 ;
        RECT 4.000 838.080 1495.600 839.480 ;
        RECT 4.000 828.600 1496.000 838.080 ;
        RECT 4.400 827.200 1496.000 828.600 ;
        RECT 4.000 823.160 1496.000 827.200 ;
        RECT 4.000 821.760 1495.600 823.160 ;
        RECT 4.000 808.880 1496.000 821.760 ;
        RECT 4.400 807.480 1496.000 808.880 ;
        RECT 4.000 806.840 1496.000 807.480 ;
        RECT 4.000 805.440 1495.600 806.840 ;
        RECT 4.000 790.520 1496.000 805.440 ;
        RECT 4.000 789.160 1495.600 790.520 ;
        RECT 4.400 789.120 1495.600 789.160 ;
        RECT 4.400 787.760 1496.000 789.120 ;
        RECT 4.000 774.200 1496.000 787.760 ;
        RECT 4.000 772.800 1495.600 774.200 ;
        RECT 4.000 770.120 1496.000 772.800 ;
        RECT 4.400 768.720 1496.000 770.120 ;
        RECT 4.000 758.560 1496.000 768.720 ;
        RECT 4.000 757.160 1495.600 758.560 ;
        RECT 4.000 750.400 1496.000 757.160 ;
        RECT 4.400 749.000 1496.000 750.400 ;
        RECT 4.000 742.240 1496.000 749.000 ;
        RECT 4.000 740.840 1495.600 742.240 ;
        RECT 4.000 731.360 1496.000 740.840 ;
        RECT 4.400 729.960 1496.000 731.360 ;
        RECT 4.000 725.920 1496.000 729.960 ;
        RECT 4.000 724.520 1495.600 725.920 ;
        RECT 4.000 711.640 1496.000 724.520 ;
        RECT 4.400 710.240 1496.000 711.640 ;
        RECT 4.000 709.600 1496.000 710.240 ;
        RECT 4.000 708.200 1495.600 709.600 ;
        RECT 4.000 693.280 1496.000 708.200 ;
        RECT 4.000 691.920 1495.600 693.280 ;
        RECT 4.400 691.880 1495.600 691.920 ;
        RECT 4.400 690.520 1496.000 691.880 ;
        RECT 4.000 676.960 1496.000 690.520 ;
        RECT 4.000 675.560 1495.600 676.960 ;
        RECT 4.000 672.880 1496.000 675.560 ;
        RECT 4.400 671.480 1496.000 672.880 ;
        RECT 4.000 660.640 1496.000 671.480 ;
        RECT 4.000 659.240 1495.600 660.640 ;
        RECT 4.000 653.160 1496.000 659.240 ;
        RECT 4.400 651.760 1496.000 653.160 ;
        RECT 4.000 644.320 1496.000 651.760 ;
        RECT 4.000 642.920 1495.600 644.320 ;
        RECT 4.000 633.440 1496.000 642.920 ;
        RECT 4.400 632.040 1496.000 633.440 ;
        RECT 4.000 628.000 1496.000 632.040 ;
        RECT 4.000 626.600 1495.600 628.000 ;
        RECT 4.000 614.400 1496.000 626.600 ;
        RECT 4.400 613.000 1496.000 614.400 ;
        RECT 4.000 611.680 1496.000 613.000 ;
        RECT 4.000 610.280 1495.600 611.680 ;
        RECT 4.000 595.360 1496.000 610.280 ;
        RECT 4.000 594.680 1495.600 595.360 ;
        RECT 4.400 593.960 1495.600 594.680 ;
        RECT 4.400 593.280 1496.000 593.960 ;
        RECT 4.000 579.040 1496.000 593.280 ;
        RECT 4.000 577.640 1495.600 579.040 ;
        RECT 4.000 574.960 1496.000 577.640 ;
        RECT 4.400 573.560 1496.000 574.960 ;
        RECT 4.000 562.720 1496.000 573.560 ;
        RECT 4.000 561.320 1495.600 562.720 ;
        RECT 4.000 555.920 1496.000 561.320 ;
        RECT 4.400 554.520 1496.000 555.920 ;
        RECT 4.000 546.400 1496.000 554.520 ;
        RECT 4.000 545.000 1495.600 546.400 ;
        RECT 4.000 536.200 1496.000 545.000 ;
        RECT 4.400 534.800 1496.000 536.200 ;
        RECT 4.000 530.080 1496.000 534.800 ;
        RECT 4.000 528.680 1495.600 530.080 ;
        RECT 4.000 516.480 1496.000 528.680 ;
        RECT 4.400 515.080 1496.000 516.480 ;
        RECT 4.000 513.760 1496.000 515.080 ;
        RECT 4.000 512.360 1495.600 513.760 ;
        RECT 4.000 497.440 1496.000 512.360 ;
        RECT 4.400 496.040 1495.600 497.440 ;
        RECT 4.000 481.120 1496.000 496.040 ;
        RECT 4.000 479.720 1495.600 481.120 ;
        RECT 4.000 477.720 1496.000 479.720 ;
        RECT 4.400 476.320 1496.000 477.720 ;
        RECT 4.000 464.800 1496.000 476.320 ;
        RECT 4.000 463.400 1495.600 464.800 ;
        RECT 4.000 458.000 1496.000 463.400 ;
        RECT 4.400 456.600 1496.000 458.000 ;
        RECT 4.000 448.480 1496.000 456.600 ;
        RECT 4.000 447.080 1495.600 448.480 ;
        RECT 4.000 438.960 1496.000 447.080 ;
        RECT 4.400 437.560 1496.000 438.960 ;
        RECT 4.000 432.160 1496.000 437.560 ;
        RECT 4.000 430.760 1495.600 432.160 ;
        RECT 4.000 419.240 1496.000 430.760 ;
        RECT 4.400 417.840 1496.000 419.240 ;
        RECT 4.000 415.840 1496.000 417.840 ;
        RECT 4.000 414.440 1495.600 415.840 ;
        RECT 4.000 399.520 1496.000 414.440 ;
        RECT 4.400 398.120 1495.600 399.520 ;
        RECT 4.000 383.200 1496.000 398.120 ;
        RECT 4.000 381.800 1495.600 383.200 ;
        RECT 4.000 380.480 1496.000 381.800 ;
        RECT 4.400 379.080 1496.000 380.480 ;
        RECT 4.000 366.880 1496.000 379.080 ;
        RECT 4.000 365.480 1495.600 366.880 ;
        RECT 4.000 360.760 1496.000 365.480 ;
        RECT 4.400 359.360 1496.000 360.760 ;
        RECT 4.000 350.560 1496.000 359.360 ;
        RECT 4.000 349.160 1495.600 350.560 ;
        RECT 4.000 341.720 1496.000 349.160 ;
        RECT 4.400 340.320 1496.000 341.720 ;
        RECT 4.000 334.240 1496.000 340.320 ;
        RECT 4.000 332.840 1495.600 334.240 ;
        RECT 4.000 322.000 1496.000 332.840 ;
        RECT 4.400 320.600 1496.000 322.000 ;
        RECT 4.000 317.920 1496.000 320.600 ;
        RECT 4.000 316.520 1495.600 317.920 ;
        RECT 4.000 302.280 1496.000 316.520 ;
        RECT 4.400 301.600 1496.000 302.280 ;
        RECT 4.400 300.880 1495.600 301.600 ;
        RECT 4.000 300.200 1495.600 300.880 ;
        RECT 4.000 285.280 1496.000 300.200 ;
        RECT 4.000 283.880 1495.600 285.280 ;
        RECT 4.000 283.240 1496.000 283.880 ;
        RECT 4.400 281.840 1496.000 283.240 ;
        RECT 4.000 268.960 1496.000 281.840 ;
        RECT 4.000 267.560 1495.600 268.960 ;
        RECT 4.000 263.520 1496.000 267.560 ;
        RECT 4.400 262.120 1496.000 263.520 ;
        RECT 4.000 252.640 1496.000 262.120 ;
        RECT 4.000 251.240 1495.600 252.640 ;
        RECT 4.000 243.800 1496.000 251.240 ;
        RECT 4.400 242.400 1496.000 243.800 ;
        RECT 4.000 236.320 1496.000 242.400 ;
        RECT 4.000 234.920 1495.600 236.320 ;
        RECT 4.000 224.760 1496.000 234.920 ;
        RECT 4.400 223.360 1496.000 224.760 ;
        RECT 4.000 220.000 1496.000 223.360 ;
        RECT 4.000 218.600 1495.600 220.000 ;
        RECT 4.000 205.040 1496.000 218.600 ;
        RECT 4.400 203.680 1496.000 205.040 ;
        RECT 4.400 203.640 1495.600 203.680 ;
        RECT 4.000 202.280 1495.600 203.640 ;
        RECT 4.000 187.360 1496.000 202.280 ;
        RECT 4.000 185.960 1495.600 187.360 ;
        RECT 4.000 185.320 1496.000 185.960 ;
        RECT 4.400 183.920 1496.000 185.320 ;
        RECT 4.000 171.040 1496.000 183.920 ;
        RECT 4.000 169.640 1495.600 171.040 ;
        RECT 4.000 166.280 1496.000 169.640 ;
        RECT 4.400 164.880 1496.000 166.280 ;
        RECT 4.000 154.720 1496.000 164.880 ;
        RECT 4.000 153.320 1495.600 154.720 ;
        RECT 4.000 146.560 1496.000 153.320 ;
        RECT 4.400 145.160 1496.000 146.560 ;
        RECT 4.000 138.400 1496.000 145.160 ;
        RECT 4.000 137.000 1495.600 138.400 ;
        RECT 4.000 126.840 1496.000 137.000 ;
        RECT 4.400 125.440 1496.000 126.840 ;
        RECT 4.000 122.080 1496.000 125.440 ;
        RECT 4.000 120.680 1495.600 122.080 ;
        RECT 4.000 107.800 1496.000 120.680 ;
        RECT 4.400 106.400 1496.000 107.800 ;
        RECT 4.000 105.760 1496.000 106.400 ;
        RECT 4.000 104.360 1495.600 105.760 ;
        RECT 4.000 89.440 1496.000 104.360 ;
        RECT 4.000 88.080 1495.600 89.440 ;
        RECT 4.400 88.040 1495.600 88.080 ;
        RECT 4.400 86.680 1496.000 88.040 ;
        RECT 4.000 73.120 1496.000 86.680 ;
        RECT 4.000 71.720 1495.600 73.120 ;
        RECT 4.000 68.360 1496.000 71.720 ;
        RECT 4.400 66.960 1496.000 68.360 ;
        RECT 4.000 56.800 1496.000 66.960 ;
        RECT 4.000 55.400 1495.600 56.800 ;
        RECT 4.000 49.320 1496.000 55.400 ;
        RECT 4.400 47.920 1496.000 49.320 ;
        RECT 4.000 40.480 1496.000 47.920 ;
        RECT 4.000 39.080 1495.600 40.480 ;
        RECT 4.000 29.600 1496.000 39.080 ;
        RECT 4.400 28.200 1496.000 29.600 ;
        RECT 4.000 24.160 1496.000 28.200 ;
        RECT 4.000 22.760 1495.600 24.160 ;
        RECT 4.000 10.560 1496.000 22.760 ;
        RECT 4.400 9.160 1496.000 10.560 ;
        RECT 4.000 8.520 1496.000 9.160 ;
        RECT 4.000 7.655 1495.600 8.520 ;
      LAYER met4 ;
        RECT 96.895 10.240 97.440 1151.065 ;
        RECT 99.840 10.240 174.240 1151.065 ;
        RECT 176.640 10.240 251.040 1151.065 ;
        RECT 253.440 10.240 327.840 1151.065 ;
        RECT 330.240 10.240 404.640 1151.065 ;
        RECT 407.040 10.240 481.440 1151.065 ;
        RECT 483.840 10.240 558.240 1151.065 ;
        RECT 560.640 10.240 635.040 1151.065 ;
        RECT 637.440 10.240 711.840 1151.065 ;
        RECT 714.240 10.240 788.640 1151.065 ;
        RECT 791.040 10.240 865.440 1151.065 ;
        RECT 867.840 10.240 942.240 1151.065 ;
        RECT 944.640 10.240 1019.040 1151.065 ;
        RECT 1021.440 10.240 1095.840 1151.065 ;
        RECT 1098.240 10.240 1158.905 1151.065 ;
        RECT 96.895 9.695 1158.905 10.240 ;
  END
END core
END LIBRARY

