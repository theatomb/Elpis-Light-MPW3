VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cache
  CLASS BLOCK ;
  FOREIGN cache ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN address_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 596.000 50.050 600.000 ;
    END
  END address_in[0]
  PIN address_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END address_in[10]
  PIN address_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END address_in[11]
  PIN address_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END address_in[12]
  PIN address_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 504.600 600.000 505.200 ;
    END
  END address_in[13]
  PIN address_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 596.000 142.050 600.000 ;
    END
  END address_in[14]
  PIN address_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 596.000 185.290 600.000 ;
    END
  END address_in[15]
  PIN address_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END address_in[16]
  PIN address_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 596.000 264.410 600.000 ;
    END
  END address_in[17]
  PIN address_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END address_in[18]
  PIN address_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END address_in[19]
  PIN address_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END address_in[1]
  PIN address_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 84.360 600.000 84.960 ;
    END
  END address_in[20]
  PIN address_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END address_in[21]
  PIN address_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END address_in[22]
  PIN address_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 596.000 334.330 600.000 ;
    END
  END address_in[23]
  PIN address_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END address_in[24]
  PIN address_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 596.000 443.810 600.000 ;
    END
  END address_in[25]
  PIN address_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END address_in[26]
  PIN address_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END address_in[27]
  PIN address_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 427.080 600.000 427.680 ;
    END
  END address_in[28]
  PIN address_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END address_in[29]
  PIN address_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END address_in[2]
  PIN address_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 518.200 600.000 518.800 ;
    END
  END address_in[30]
  PIN address_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 596.000 132.850 600.000 ;
    END
  END address_in[31]
  PIN address_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END address_in[3]
  PIN address_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END address_in[4]
  PIN address_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 232.600 600.000 233.200 ;
    END
  END address_in[5]
  PIN address_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END address_in[6]
  PIN address_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END address_in[7]
  PIN address_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 6.840 600.000 7.440 ;
    END
  END address_in[8]
  PIN address_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 342.760 600.000 343.360 ;
    END
  END address_in[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 596.000 365.610 600.000 ;
    END
  END clk
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 110.200 600.000 110.800 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 596.000 589.170 600.000 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 596.000 553.290 600.000 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 201.320 600.000 201.920 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 19.080 600.000 19.680 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 576.680 600.000 577.280 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 478.760 600.000 479.360 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 596.000 461.290 600.000 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 596.000 575.370 600.000 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 596.000 453.010 600.000 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 596.000 89.610 600.000 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 25.880 600.000 26.480 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 596.000 567.090 600.000 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 596.000 110.770 600.000 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 596.000 256.130 600.000 ;
    END
  END data_in[31]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 122.440 600.000 123.040 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 96.600 600.000 97.200 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 596.000 5.890 600.000 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END data_in[9]
  PIN exc_protected_page_tlb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 142.840 600.000 143.440 ;
    END
  END exc_protected_page_tlb
  PIN hit_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 213.560 600.000 214.160 ;
    END
  END hit_out
  PIN hit_tlb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 596.000 129.170 600.000 ;
    END
  END hit_tlb
  PIN is_byte
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END is_byte
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 596.000 150.330 600.000 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 595.720 600.000 596.320 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 129.240 600.000 129.840 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 356.360 600.000 356.960 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 596.000 15.090 600.000 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 596.000 330.650 600.000 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 258.440 600.000 259.040 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 596.000 277.290 600.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 596.000 107.090 600.000 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 596.000 1.290 600.000 ;
    END
  END mem_addr_out[9]
  PIN mem_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 596.000 408.850 600.000 ;
    END
  END mem_data_in[0]
  PIN mem_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END mem_data_in[100]
  PIN mem_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 596.000 216.570 600.000 ;
    END
  END mem_data_in[101]
  PIN mem_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 596.000 413.450 600.000 ;
    END
  END mem_data_in[102]
  PIN mem_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END mem_data_in[103]
  PIN mem_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 65.320 600.000 65.920 ;
    END
  END mem_data_in[104]
  PIN mem_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END mem_data_in[105]
  PIN mem_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 304.680 600.000 305.280 ;
    END
  END mem_data_in[106]
  PIN mem_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 596.000 23.370 600.000 ;
    END
  END mem_data_in[107]
  PIN mem_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 32.680 600.000 33.280 ;
    END
  END mem_data_in[108]
  PIN mem_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END mem_data_in[109]
  PIN mem_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END mem_data_in[10]
  PIN mem_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END mem_data_in[110]
  PIN mem_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 596.000 181.610 600.000 ;
    END
  END mem_data_in[111]
  PIN mem_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 596.000 54.650 600.000 ;
    END
  END mem_data_in[112]
  PIN mem_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END mem_data_in[113]
  PIN mem_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END mem_data_in[114]
  PIN mem_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END mem_data_in[115]
  PIN mem_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 187.720 600.000 188.320 ;
    END
  END mem_data_in[116]
  PIN mem_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END mem_data_in[117]
  PIN mem_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 596.000 435.530 600.000 ;
    END
  END mem_data_in[118]
  PIN mem_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END mem_data_in[119]
  PIN mem_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 596.000 251.530 600.000 ;
    END
  END mem_data_in[11]
  PIN mem_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END mem_data_in[120]
  PIN mem_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 596.000 62.930 600.000 ;
    END
  END mem_data_in[121]
  PIN mem_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END mem_data_in[122]
  PIN mem_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 596.000 522.930 600.000 ;
    END
  END mem_data_in[123]
  PIN mem_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 421.640 600.000 422.240 ;
    END
  END mem_data_in[124]
  PIN mem_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END mem_data_in[125]
  PIN mem_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 596.000 75.810 600.000 ;
    END
  END mem_data_in[126]
  PIN mem_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END mem_data_in[127]
  PIN mem_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 596.000 532.130 600.000 ;
    END
  END mem_data_in[12]
  PIN mem_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 596.000 510.050 600.000 ;
    END
  END mem_data_in[13]
  PIN mem_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 155.080 600.000 155.680 ;
    END
  END mem_data_in[14]
  PIN mem_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 596.000 295.690 600.000 ;
    END
  END mem_data_in[15]
  PIN mem_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 492.360 600.000 492.960 ;
    END
  END mem_data_in[16]
  PIN mem_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 0.040 600.000 0.640 ;
    END
  END mem_data_in[17]
  PIN mem_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END mem_data_in[18]
  PIN mem_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END mem_data_in[19]
  PIN mem_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 596.000 124.570 600.000 ;
    END
  END mem_data_in[1]
  PIN mem_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END mem_data_in[20]
  PIN mem_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END mem_data_in[21]
  PIN mem_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 596.000 383.090 600.000 ;
    END
  END mem_data_in[22]
  PIN mem_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 596.000 246.930 600.000 ;
    END
  END mem_data_in[23]
  PIN mem_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 596.000 557.890 600.000 ;
    END
  END mem_data_in[24]
  PIN mem_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END mem_data_in[25]
  PIN mem_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 596.000 313.170 600.000 ;
    END
  END mem_data_in[26]
  PIN mem_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END mem_data_in[27]
  PIN mem_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END mem_data_in[28]
  PIN mem_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END mem_data_in[29]
  PIN mem_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END mem_data_in[2]
  PIN mem_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 596.000 164.130 600.000 ;
    END
  END mem_data_in[30]
  PIN mem_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 596.000 514.650 600.000 ;
    END
  END mem_data_in[31]
  PIN mem_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 414.840 600.000 415.440 ;
    END
  END mem_data_in[32]
  PIN mem_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 596.000 189.890 600.000 ;
    END
  END mem_data_in[33]
  PIN mem_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 596.000 115.370 600.000 ;
    END
  END mem_data_in[34]
  PIN mem_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 596.000 361.010 600.000 ;
    END
  END mem_data_in[35]
  PIN mem_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END mem_data_in[36]
  PIN mem_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 239.400 600.000 240.000 ;
    END
  END mem_data_in[37]
  PIN mem_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END mem_data_in[38]
  PIN mem_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 175.480 600.000 176.080 ;
    END
  END mem_data_in[39]
  PIN mem_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END mem_data_in[3]
  PIN mem_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 499.160 600.000 499.760 ;
    END
  END mem_data_in[40]
  PIN mem_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 297.880 600.000 298.480 ;
    END
  END mem_data_in[41]
  PIN mem_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END mem_data_in[42]
  PIN mem_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 596.000 273.610 600.000 ;
    END
  END mem_data_in[43]
  PIN mem_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 550.840 600.000 551.440 ;
    END
  END mem_data_in[44]
  PIN mem_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END mem_data_in[45]
  PIN mem_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END mem_data_in[46]
  PIN mem_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 44.920 600.000 45.520 ;
    END
  END mem_data_in[47]
  PIN mem_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END mem_data_in[48]
  PIN mem_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END mem_data_in[49]
  PIN mem_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 596.000 37.170 600.000 ;
    END
  END mem_data_in[4]
  PIN mem_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 596.000 299.370 600.000 ;
    END
  END mem_data_in[50]
  PIN mem_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 596.000 97.890 600.000 ;
    END
  END mem_data_in[51]
  PIN mem_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END mem_data_in[52]
  PIN mem_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 161.880 600.000 162.480 ;
    END
  END mem_data_in[53]
  PIN mem_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 596.000 211.970 600.000 ;
    END
  END mem_data_in[54]
  PIN mem_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END mem_data_in[55]
  PIN mem_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END mem_data_in[56]
  PIN mem_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 447.480 600.000 448.080 ;
    END
  END mem_data_in[57]
  PIN mem_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 473.320 600.000 473.920 ;
    END
  END mem_data_in[58]
  PIN mem_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END mem_data_in[59]
  PIN mem_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 596.000 338.930 600.000 ;
    END
  END mem_data_in[5]
  PIN mem_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END mem_data_in[60]
  PIN mem_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END mem_data_in[61]
  PIN mem_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END mem_data_in[62]
  PIN mem_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END mem_data_in[63]
  PIN mem_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 544.040 600.000 544.640 ;
    END
  END mem_data_in[64]
  PIN mem_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 227.160 600.000 227.760 ;
    END
  END mem_data_in[65]
  PIN mem_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END mem_data_in[66]
  PIN mem_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 596.000 369.290 600.000 ;
    END
  END mem_data_in[67]
  PIN mem_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 596.000 32.570 600.000 ;
    END
  END mem_data_in[68]
  PIN mem_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 596.000 27.970 600.000 ;
    END
  END mem_data_in[69]
  PIN mem_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END mem_data_in[6]
  PIN mem_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END mem_data_in[70]
  PIN mem_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END mem_data_in[71]
  PIN mem_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 596.000 316.850 600.000 ;
    END
  END mem_data_in[72]
  PIN mem_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 563.080 600.000 563.680 ;
    END
  END mem_data_in[73]
  PIN mem_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END mem_data_in[74]
  PIN mem_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END mem_data_in[75]
  PIN mem_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 278.840 600.000 279.440 ;
    END
  END mem_data_in[76]
  PIN mem_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 596.000 67.530 600.000 ;
    END
  END mem_data_in[77]
  PIN mem_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END mem_data_in[78]
  PIN mem_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END mem_data_in[79]
  PIN mem_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 485.560 600.000 486.160 ;
    END
  END mem_data_in[7]
  PIN mem_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 596.000 207.370 600.000 ;
    END
  END mem_data_in[80]
  PIN mem_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END mem_data_in[81]
  PIN mem_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END mem_data_in[82]
  PIN mem_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END mem_data_in[83]
  PIN mem_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END mem_data_in[84]
  PIN mem_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END mem_data_in[85]
  PIN mem_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 596.000 387.690 600.000 ;
    END
  END mem_data_in[86]
  PIN mem_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END mem_data_in[87]
  PIN mem_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 596.000 518.330 600.000 ;
    END
  END mem_data_in[88]
  PIN mem_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 596.000 400.570 600.000 ;
    END
  END mem_data_in[89]
  PIN mem_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END mem_data_in[8]
  PIN mem_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 596.000 356.410 600.000 ;
    END
  END mem_data_in[90]
  PIN mem_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END mem_data_in[91]
  PIN mem_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END mem_data_in[92]
  PIN mem_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END mem_data_in[93]
  PIN mem_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END mem_data_in[94]
  PIN mem_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END mem_data_in[95]
  PIN mem_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END mem_data_in[96]
  PIN mem_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 511.400 600.000 512.000 ;
    END
  END mem_data_in[97]
  PIN mem_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 596.000 479.690 600.000 ;
    END
  END mem_data_in[98]
  PIN mem_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END mem_data_in[99]
  PIN mem_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 368.600 600.000 369.200 ;
    END
  END mem_data_in[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 253.000 600.000 253.600 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 596.000 40.850 600.000 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 596.000 549.610 600.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 596.000 343.530 600.000 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 596.000 259.810 600.000 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 401.240 600.000 401.840 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 596.000 194.490 600.000 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 596.000 584.570 600.000 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 330.520 600.000 331.120 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 58.520 600.000 59.120 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 525.000 600.000 525.600 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 452.920 600.000 453.520 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 180.920 600.000 181.520 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 596.000 303.970 600.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 596.000 326.050 600.000 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 588.920 600.000 589.520 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 596.000 308.570 600.000 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 596.000 430.930 600.000 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 596.000 242.330 600.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 596.000 291.090 600.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 583.480 600.000 584.080 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 246.200 600.000 246.800 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 39.480 600.000 40.080 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 168.680 600.000 169.280 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 596.000 592.850 600.000 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 596.000 321.450 600.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 596.000 85.010 600.000 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 596.000 378.490 600.000 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 103.400 600.000 104.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 596.000 45.450 600.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 596.000 579.970 600.000 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 596.000 93.290 600.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 136.040 600.000 136.640 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 596.000 505.450 600.000 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 596.000 137.450 600.000 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 206.760 600.000 207.360 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 596.000 72.130 600.000 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 349.560 600.000 350.160 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 363.160 600.000 363.760 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 596.000 172.410 600.000 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 596.000 281.890 600.000 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 596.000 269.010 600.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 596.000 497.170 600.000 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 596.000 475.090 600.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 596.000 405.170 600.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 382.200 600.000 382.800 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 596.000 373.890 600.000 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 311.480 600.000 312.080 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 596.000 571.690 600.000 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 596.000 540.410 600.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 569.880 600.000 570.480 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 596.000 154.930 600.000 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 596.000 487.970 600.000 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 596.000 159.530 600.000 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 596.000 527.530 600.000 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 596.000 221.170 600.000 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 596.000 202.770 600.000 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 375.400 600.000 376.000 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 285.640 600.000 286.240 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 596.000 348.130 600.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 596.000 167.810 600.000 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 272.040 600.000 272.640 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END mem_data_out[9]
  PIN mem_ready_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 389.000 600.000 389.600 ;
    END
  END mem_ready_in
  PIN mem_we_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END mem_we_out
  PIN physical_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END physical_addr_in[0]
  PIN physical_addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END physical_addr_in[10]
  PIN physical_addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 596.000 492.570 600.000 ;
    END
  END physical_addr_in[11]
  PIN physical_addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 466.520 600.000 467.120 ;
    END
  END physical_addr_in[12]
  PIN physical_addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 596.000 177.010 600.000 ;
    END
  END physical_addr_in[13]
  PIN physical_addr_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 596.000 224.850 600.000 ;
    END
  END physical_addr_in[14]
  PIN physical_addr_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 12.280 600.000 12.880 ;
    END
  END physical_addr_in[15]
  PIN physical_addr_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END physical_addr_in[16]
  PIN physical_addr_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 149.640 600.000 150.240 ;
    END
  END physical_addr_in[17]
  PIN physical_addr_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 596.000 395.970 600.000 ;
    END
  END physical_addr_in[18]
  PIN physical_addr_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 596.000 286.490 600.000 ;
    END
  END physical_addr_in[19]
  PIN physical_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 596.000 80.410 600.000 ;
    END
  END physical_addr_in[1]
  PIN physical_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END physical_addr_in[2]
  PIN physical_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END physical_addr_in[3]
  PIN physical_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 440.680 600.000 441.280 ;
    END
  END physical_addr_in[4]
  PIN physical_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 394.440 600.000 395.040 ;
    END
  END physical_addr_in[5]
  PIN physical_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END physical_addr_in[6]
  PIN physical_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 337.320 600.000 337.920 ;
    END
  END physical_addr_in[7]
  PIN physical_addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END physical_addr_in[8]
  PIN physical_addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 4.000 ;
    END
  END physical_addr_in[9]
  PIN physical_addr_write_tlb_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 596.000 391.370 600.000 ;
    END
  END physical_addr_write_tlb_in[0]
  PIN physical_addr_write_tlb_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 596.000 535.810 600.000 ;
    END
  END physical_addr_write_tlb_in[10]
  PIN physical_addr_write_tlb_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END physical_addr_write_tlb_in[11]
  PIN physical_addr_write_tlb_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END physical_addr_write_tlb_in[12]
  PIN physical_addr_write_tlb_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 51.720 600.000 52.320 ;
    END
  END physical_addr_write_tlb_in[13]
  PIN physical_addr_write_tlb_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 596.000 119.970 600.000 ;
    END
  END physical_addr_write_tlb_in[14]
  PIN physical_addr_write_tlb_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END physical_addr_write_tlb_in[15]
  PIN physical_addr_write_tlb_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END physical_addr_write_tlb_in[16]
  PIN physical_addr_write_tlb_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 596.000 234.050 600.000 ;
    END
  END physical_addr_write_tlb_in[17]
  PIN physical_addr_write_tlb_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 316.920 600.000 317.520 ;
    END
  END physical_addr_write_tlb_in[18]
  PIN physical_addr_write_tlb_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 596.000 597.450 600.000 ;
    END
  END physical_addr_write_tlb_in[19]
  PIN physical_addr_write_tlb_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END physical_addr_write_tlb_in[1]
  PIN physical_addr_write_tlb_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 596.000 470.490 600.000 ;
    END
  END physical_addr_write_tlb_in[2]
  PIN physical_addr_write_tlb_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END physical_addr_write_tlb_in[3]
  PIN physical_addr_write_tlb_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END physical_addr_write_tlb_in[4]
  PIN physical_addr_write_tlb_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 596.000 457.610 600.000 ;
    END
  END physical_addr_write_tlb_in[5]
  PIN physical_addr_write_tlb_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END physical_addr_write_tlb_in[6]
  PIN physical_addr_write_tlb_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END physical_addr_write_tlb_in[7]
  PIN physical_addr_write_tlb_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END physical_addr_write_tlb_in[8]
  PIN physical_addr_write_tlb_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END physical_addr_write_tlb_in[9]
  PIN privilege_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 77.560 600.000 78.160 ;
    END
  END privilege_mode
  PIN read_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END read_data_out[0]
  PIN read_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 530.440 600.000 531.040 ;
    END
  END read_data_out[10]
  PIN read_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END read_data_out[11]
  PIN read_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END read_data_out[12]
  PIN read_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END read_data_out[13]
  PIN read_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END read_data_out[14]
  PIN read_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END read_data_out[15]
  PIN read_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 265.240 600.000 265.840 ;
    END
  END read_data_out[16]
  PIN read_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END read_data_out[17]
  PIN read_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 596.000 422.650 600.000 ;
    END
  END read_data_out[18]
  PIN read_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 596.000 545.010 600.000 ;
    END
  END read_data_out[19]
  PIN read_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 596.000 102.490 600.000 ;
    END
  END read_data_out[1]
  PIN read_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END read_data_out[20]
  PIN read_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END read_data_out[21]
  PIN read_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 596.000 562.490 600.000 ;
    END
  END read_data_out[22]
  PIN read_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END read_data_out[23]
  PIN read_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 459.720 600.000 460.320 ;
    END
  END read_data_out[24]
  PIN read_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 117.000 600.000 117.600 ;
    END
  END read_data_out[25]
  PIN read_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END read_data_out[26]
  PIN read_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 596.000 500.850 600.000 ;
    END
  END read_data_out[27]
  PIN read_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 596.000 199.090 600.000 ;
    END
  END read_data_out[28]
  PIN read_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END read_data_out[29]
  PIN read_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 323.720 600.000 324.320 ;
    END
  END read_data_out[2]
  PIN read_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END read_data_out[30]
  PIN read_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 91.160 600.000 91.760 ;
    END
  END read_data_out[31]
  PIN read_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END read_data_out[3]
  PIN read_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END read_data_out[4]
  PIN read_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END read_data_out[5]
  PIN read_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END read_data_out[6]
  PIN read_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 194.520 600.000 195.120 ;
    END
  END read_data_out[7]
  PIN read_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 596.000 483.370 600.000 ;
    END
  END read_data_out[8]
  PIN read_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 537.240 600.000 537.840 ;
    END
  END read_data_out[9]
  PIN read_enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END read_enable_in
  PIN req_mem
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END req_mem
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 291.080 600.000 291.680 ;
    END
  END reset
  PIN reset_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END reset_mem_req
  PIN tlb_re
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 557.640 600.000 558.240 ;
    END
  END tlb_re
  PIN tlb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 596.000 465.890 600.000 ;
    END
  END tlb_we
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN virtual_addr_write_tlb_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END virtual_addr_write_tlb_in[0]
  PIN virtual_addr_write_tlb_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 596.000 448.410 600.000 ;
    END
  END virtual_addr_write_tlb_in[10]
  PIN virtual_addr_write_tlb_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END virtual_addr_write_tlb_in[11]
  PIN virtual_addr_write_tlb_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END virtual_addr_write_tlb_in[12]
  PIN virtual_addr_write_tlb_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END virtual_addr_write_tlb_in[13]
  PIN virtual_addr_write_tlb_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END virtual_addr_write_tlb_in[14]
  PIN virtual_addr_write_tlb_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END virtual_addr_write_tlb_in[15]
  PIN virtual_addr_write_tlb_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END virtual_addr_write_tlb_in[16]
  PIN virtual_addr_write_tlb_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 596.000 18.770 600.000 ;
    END
  END virtual_addr_write_tlb_in[17]
  PIN virtual_addr_write_tlb_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 596.000 229.450 600.000 ;
    END
  END virtual_addr_write_tlb_in[18]
  PIN virtual_addr_write_tlb_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END virtual_addr_write_tlb_in[19]
  PIN virtual_addr_write_tlb_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END virtual_addr_write_tlb_in[1]
  PIN virtual_addr_write_tlb_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END virtual_addr_write_tlb_in[20]
  PIN virtual_addr_write_tlb_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 596.000 351.810 600.000 ;
    END
  END virtual_addr_write_tlb_in[21]
  PIN virtual_addr_write_tlb_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 596.000 238.650 600.000 ;
    END
  END virtual_addr_write_tlb_in[22]
  PIN virtual_addr_write_tlb_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END virtual_addr_write_tlb_in[23]
  PIN virtual_addr_write_tlb_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 596.000 440.130 600.000 ;
    END
  END virtual_addr_write_tlb_in[24]
  PIN virtual_addr_write_tlb_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 70.760 600.000 71.360 ;
    END
  END virtual_addr_write_tlb_in[25]
  PIN virtual_addr_write_tlb_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END virtual_addr_write_tlb_in[26]
  PIN virtual_addr_write_tlb_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 433.880 600.000 434.480 ;
    END
  END virtual_addr_write_tlb_in[27]
  PIN virtual_addr_write_tlb_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END virtual_addr_write_tlb_in[28]
  PIN virtual_addr_write_tlb_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END virtual_addr_write_tlb_in[29]
  PIN virtual_addr_write_tlb_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END virtual_addr_write_tlb_in[2]
  PIN virtual_addr_write_tlb_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 408.040 600.000 408.640 ;
    END
  END virtual_addr_write_tlb_in[30]
  PIN virtual_addr_write_tlb_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END virtual_addr_write_tlb_in[31]
  PIN virtual_addr_write_tlb_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 596.000 426.330 600.000 ;
    END
  END virtual_addr_write_tlb_in[3]
  PIN virtual_addr_write_tlb_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 596.000 418.050 600.000 ;
    END
  END virtual_addr_write_tlb_in[4]
  PIN virtual_addr_write_tlb_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 596.000 58.330 600.000 ;
    END
  END virtual_addr_write_tlb_in[5]
  PIN virtual_addr_write_tlb_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 596.000 146.650 600.000 ;
    END
  END virtual_addr_write_tlb_in[6]
  PIN virtual_addr_write_tlb_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END virtual_addr_write_tlb_in[7]
  PIN virtual_addr_write_tlb_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END virtual_addr_write_tlb_in[8]
  PIN virtual_addr_write_tlb_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 596.000 10.490 600.000 ;
    END
  END virtual_addr_write_tlb_in[9]
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN write_enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 220.360 600.000 220.960 ;
    END
  END write_enable_in
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 596.935 595.935 ;
      LAYER met1 ;
        RECT 0.990 6.840 596.995 595.980 ;
      LAYER met2 ;
        RECT 1.570 595.720 5.330 596.205 ;
        RECT 6.170 595.720 9.930 596.205 ;
        RECT 10.770 595.720 14.530 596.205 ;
        RECT 15.370 595.720 18.210 596.205 ;
        RECT 19.050 595.720 22.810 596.205 ;
        RECT 23.650 595.720 27.410 596.205 ;
        RECT 28.250 595.720 32.010 596.205 ;
        RECT 32.850 595.720 36.610 596.205 ;
        RECT 37.450 595.720 40.290 596.205 ;
        RECT 41.130 595.720 44.890 596.205 ;
        RECT 45.730 595.720 49.490 596.205 ;
        RECT 50.330 595.720 54.090 596.205 ;
        RECT 54.930 595.720 57.770 596.205 ;
        RECT 58.610 595.720 62.370 596.205 ;
        RECT 63.210 595.720 66.970 596.205 ;
        RECT 67.810 595.720 71.570 596.205 ;
        RECT 72.410 595.720 75.250 596.205 ;
        RECT 76.090 595.720 79.850 596.205 ;
        RECT 80.690 595.720 84.450 596.205 ;
        RECT 85.290 595.720 89.050 596.205 ;
        RECT 89.890 595.720 92.730 596.205 ;
        RECT 93.570 595.720 97.330 596.205 ;
        RECT 98.170 595.720 101.930 596.205 ;
        RECT 102.770 595.720 106.530 596.205 ;
        RECT 107.370 595.720 110.210 596.205 ;
        RECT 111.050 595.720 114.810 596.205 ;
        RECT 115.650 595.720 119.410 596.205 ;
        RECT 120.250 595.720 124.010 596.205 ;
        RECT 124.850 595.720 128.610 596.205 ;
        RECT 129.450 595.720 132.290 596.205 ;
        RECT 133.130 595.720 136.890 596.205 ;
        RECT 137.730 595.720 141.490 596.205 ;
        RECT 142.330 595.720 146.090 596.205 ;
        RECT 146.930 595.720 149.770 596.205 ;
        RECT 150.610 595.720 154.370 596.205 ;
        RECT 155.210 595.720 158.970 596.205 ;
        RECT 159.810 595.720 163.570 596.205 ;
        RECT 164.410 595.720 167.250 596.205 ;
        RECT 168.090 595.720 171.850 596.205 ;
        RECT 172.690 595.720 176.450 596.205 ;
        RECT 177.290 595.720 181.050 596.205 ;
        RECT 181.890 595.720 184.730 596.205 ;
        RECT 185.570 595.720 189.330 596.205 ;
        RECT 190.170 595.720 193.930 596.205 ;
        RECT 194.770 595.720 198.530 596.205 ;
        RECT 199.370 595.720 202.210 596.205 ;
        RECT 203.050 595.720 206.810 596.205 ;
        RECT 207.650 595.720 211.410 596.205 ;
        RECT 212.250 595.720 216.010 596.205 ;
        RECT 216.850 595.720 220.610 596.205 ;
        RECT 221.450 595.720 224.290 596.205 ;
        RECT 225.130 595.720 228.890 596.205 ;
        RECT 229.730 595.720 233.490 596.205 ;
        RECT 234.330 595.720 238.090 596.205 ;
        RECT 238.930 595.720 241.770 596.205 ;
        RECT 242.610 595.720 246.370 596.205 ;
        RECT 247.210 595.720 250.970 596.205 ;
        RECT 251.810 595.720 255.570 596.205 ;
        RECT 256.410 595.720 259.250 596.205 ;
        RECT 260.090 595.720 263.850 596.205 ;
        RECT 264.690 595.720 268.450 596.205 ;
        RECT 269.290 595.720 273.050 596.205 ;
        RECT 273.890 595.720 276.730 596.205 ;
        RECT 277.570 595.720 281.330 596.205 ;
        RECT 282.170 595.720 285.930 596.205 ;
        RECT 286.770 595.720 290.530 596.205 ;
        RECT 291.370 595.720 295.130 596.205 ;
        RECT 295.970 595.720 298.810 596.205 ;
        RECT 299.650 595.720 303.410 596.205 ;
        RECT 304.250 595.720 308.010 596.205 ;
        RECT 308.850 595.720 312.610 596.205 ;
        RECT 313.450 595.720 316.290 596.205 ;
        RECT 317.130 595.720 320.890 596.205 ;
        RECT 321.730 595.720 325.490 596.205 ;
        RECT 326.330 595.720 330.090 596.205 ;
        RECT 330.930 595.720 333.770 596.205 ;
        RECT 334.610 595.720 338.370 596.205 ;
        RECT 339.210 595.720 342.970 596.205 ;
        RECT 343.810 595.720 347.570 596.205 ;
        RECT 348.410 595.720 351.250 596.205 ;
        RECT 352.090 595.720 355.850 596.205 ;
        RECT 356.690 595.720 360.450 596.205 ;
        RECT 361.290 595.720 365.050 596.205 ;
        RECT 365.890 595.720 368.730 596.205 ;
        RECT 369.570 595.720 373.330 596.205 ;
        RECT 374.170 595.720 377.930 596.205 ;
        RECT 378.770 595.720 382.530 596.205 ;
        RECT 383.370 595.720 387.130 596.205 ;
        RECT 387.970 595.720 390.810 596.205 ;
        RECT 391.650 595.720 395.410 596.205 ;
        RECT 396.250 595.720 400.010 596.205 ;
        RECT 400.850 595.720 404.610 596.205 ;
        RECT 405.450 595.720 408.290 596.205 ;
        RECT 409.130 595.720 412.890 596.205 ;
        RECT 413.730 595.720 417.490 596.205 ;
        RECT 418.330 595.720 422.090 596.205 ;
        RECT 422.930 595.720 425.770 596.205 ;
        RECT 426.610 595.720 430.370 596.205 ;
        RECT 431.210 595.720 434.970 596.205 ;
        RECT 435.810 595.720 439.570 596.205 ;
        RECT 440.410 595.720 443.250 596.205 ;
        RECT 444.090 595.720 447.850 596.205 ;
        RECT 448.690 595.720 452.450 596.205 ;
        RECT 453.290 595.720 457.050 596.205 ;
        RECT 457.890 595.720 460.730 596.205 ;
        RECT 461.570 595.720 465.330 596.205 ;
        RECT 466.170 595.720 469.930 596.205 ;
        RECT 470.770 595.720 474.530 596.205 ;
        RECT 475.370 595.720 479.130 596.205 ;
        RECT 479.970 595.720 482.810 596.205 ;
        RECT 483.650 595.720 487.410 596.205 ;
        RECT 488.250 595.720 492.010 596.205 ;
        RECT 492.850 595.720 496.610 596.205 ;
        RECT 497.450 595.720 500.290 596.205 ;
        RECT 501.130 595.720 504.890 596.205 ;
        RECT 505.730 595.720 509.490 596.205 ;
        RECT 510.330 595.720 514.090 596.205 ;
        RECT 514.930 595.720 517.770 596.205 ;
        RECT 518.610 595.720 522.370 596.205 ;
        RECT 523.210 595.720 526.970 596.205 ;
        RECT 527.810 595.720 531.570 596.205 ;
        RECT 532.410 595.720 535.250 596.205 ;
        RECT 536.090 595.720 539.850 596.205 ;
        RECT 540.690 595.720 544.450 596.205 ;
        RECT 545.290 595.720 549.050 596.205 ;
        RECT 549.890 595.720 552.730 596.205 ;
        RECT 553.570 595.720 557.330 596.205 ;
        RECT 558.170 595.720 561.930 596.205 ;
        RECT 562.770 595.720 566.530 596.205 ;
        RECT 567.370 595.720 571.130 596.205 ;
        RECT 571.970 595.720 574.810 596.205 ;
        RECT 575.650 595.720 579.410 596.205 ;
        RECT 580.250 595.720 584.010 596.205 ;
        RECT 584.850 595.720 588.610 596.205 ;
        RECT 589.450 595.720 592.290 596.205 ;
        RECT 593.130 595.720 595.610 596.205 ;
        RECT 1.020 4.280 595.610 595.720 ;
        RECT 1.020 0.155 3.490 4.280 ;
        RECT 4.330 0.155 8.090 4.280 ;
        RECT 8.930 0.155 12.690 4.280 ;
        RECT 13.530 0.155 17.290 4.280 ;
        RECT 18.130 0.155 20.970 4.280 ;
        RECT 21.810 0.155 25.570 4.280 ;
        RECT 26.410 0.155 30.170 4.280 ;
        RECT 31.010 0.155 34.770 4.280 ;
        RECT 35.610 0.155 38.450 4.280 ;
        RECT 39.290 0.155 43.050 4.280 ;
        RECT 43.890 0.155 47.650 4.280 ;
        RECT 48.490 0.155 52.250 4.280 ;
        RECT 53.090 0.155 55.930 4.280 ;
        RECT 56.770 0.155 60.530 4.280 ;
        RECT 61.370 0.155 65.130 4.280 ;
        RECT 65.970 0.155 69.730 4.280 ;
        RECT 70.570 0.155 73.410 4.280 ;
        RECT 74.250 0.155 78.010 4.280 ;
        RECT 78.850 0.155 82.610 4.280 ;
        RECT 83.450 0.155 87.210 4.280 ;
        RECT 88.050 0.155 91.810 4.280 ;
        RECT 92.650 0.155 95.490 4.280 ;
        RECT 96.330 0.155 100.090 4.280 ;
        RECT 100.930 0.155 104.690 4.280 ;
        RECT 105.530 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.970 4.280 ;
        RECT 113.810 0.155 117.570 4.280 ;
        RECT 118.410 0.155 122.170 4.280 ;
        RECT 123.010 0.155 126.770 4.280 ;
        RECT 127.610 0.155 130.450 4.280 ;
        RECT 131.290 0.155 135.050 4.280 ;
        RECT 135.890 0.155 139.650 4.280 ;
        RECT 140.490 0.155 144.250 4.280 ;
        RECT 145.090 0.155 147.930 4.280 ;
        RECT 148.770 0.155 152.530 4.280 ;
        RECT 153.370 0.155 157.130 4.280 ;
        RECT 157.970 0.155 161.730 4.280 ;
        RECT 162.570 0.155 165.410 4.280 ;
        RECT 166.250 0.155 170.010 4.280 ;
        RECT 170.850 0.155 174.610 4.280 ;
        RECT 175.450 0.155 179.210 4.280 ;
        RECT 180.050 0.155 183.810 4.280 ;
        RECT 184.650 0.155 187.490 4.280 ;
        RECT 188.330 0.155 192.090 4.280 ;
        RECT 192.930 0.155 196.690 4.280 ;
        RECT 197.530 0.155 201.290 4.280 ;
        RECT 202.130 0.155 204.970 4.280 ;
        RECT 205.810 0.155 209.570 4.280 ;
        RECT 210.410 0.155 214.170 4.280 ;
        RECT 215.010 0.155 218.770 4.280 ;
        RECT 219.610 0.155 222.450 4.280 ;
        RECT 223.290 0.155 227.050 4.280 ;
        RECT 227.890 0.155 231.650 4.280 ;
        RECT 232.490 0.155 236.250 4.280 ;
        RECT 237.090 0.155 239.930 4.280 ;
        RECT 240.770 0.155 244.530 4.280 ;
        RECT 245.370 0.155 249.130 4.280 ;
        RECT 249.970 0.155 253.730 4.280 ;
        RECT 254.570 0.155 257.410 4.280 ;
        RECT 258.250 0.155 262.010 4.280 ;
        RECT 262.850 0.155 266.610 4.280 ;
        RECT 267.450 0.155 271.210 4.280 ;
        RECT 272.050 0.155 275.810 4.280 ;
        RECT 276.650 0.155 279.490 4.280 ;
        RECT 280.330 0.155 284.090 4.280 ;
        RECT 284.930 0.155 288.690 4.280 ;
        RECT 289.530 0.155 293.290 4.280 ;
        RECT 294.130 0.155 296.970 4.280 ;
        RECT 297.810 0.155 301.570 4.280 ;
        RECT 302.410 0.155 306.170 4.280 ;
        RECT 307.010 0.155 310.770 4.280 ;
        RECT 311.610 0.155 314.450 4.280 ;
        RECT 315.290 0.155 319.050 4.280 ;
        RECT 319.890 0.155 323.650 4.280 ;
        RECT 324.490 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.930 4.280 ;
        RECT 332.770 0.155 336.530 4.280 ;
        RECT 337.370 0.155 341.130 4.280 ;
        RECT 341.970 0.155 345.730 4.280 ;
        RECT 346.570 0.155 350.330 4.280 ;
        RECT 351.170 0.155 354.010 4.280 ;
        RECT 354.850 0.155 358.610 4.280 ;
        RECT 359.450 0.155 363.210 4.280 ;
        RECT 364.050 0.155 367.810 4.280 ;
        RECT 368.650 0.155 371.490 4.280 ;
        RECT 372.330 0.155 376.090 4.280 ;
        RECT 376.930 0.155 380.690 4.280 ;
        RECT 381.530 0.155 385.290 4.280 ;
        RECT 386.130 0.155 388.970 4.280 ;
        RECT 389.810 0.155 393.570 4.280 ;
        RECT 394.410 0.155 398.170 4.280 ;
        RECT 399.010 0.155 402.770 4.280 ;
        RECT 403.610 0.155 406.450 4.280 ;
        RECT 407.290 0.155 411.050 4.280 ;
        RECT 411.890 0.155 415.650 4.280 ;
        RECT 416.490 0.155 420.250 4.280 ;
        RECT 421.090 0.155 423.930 4.280 ;
        RECT 424.770 0.155 428.530 4.280 ;
        RECT 429.370 0.155 433.130 4.280 ;
        RECT 433.970 0.155 437.730 4.280 ;
        RECT 438.570 0.155 442.330 4.280 ;
        RECT 443.170 0.155 446.010 4.280 ;
        RECT 446.850 0.155 450.610 4.280 ;
        RECT 451.450 0.155 455.210 4.280 ;
        RECT 456.050 0.155 459.810 4.280 ;
        RECT 460.650 0.155 463.490 4.280 ;
        RECT 464.330 0.155 468.090 4.280 ;
        RECT 468.930 0.155 472.690 4.280 ;
        RECT 473.530 0.155 477.290 4.280 ;
        RECT 478.130 0.155 480.970 4.280 ;
        RECT 481.810 0.155 485.570 4.280 ;
        RECT 486.410 0.155 490.170 4.280 ;
        RECT 491.010 0.155 494.770 4.280 ;
        RECT 495.610 0.155 498.450 4.280 ;
        RECT 499.290 0.155 503.050 4.280 ;
        RECT 503.890 0.155 507.650 4.280 ;
        RECT 508.490 0.155 512.250 4.280 ;
        RECT 513.090 0.155 515.930 4.280 ;
        RECT 516.770 0.155 520.530 4.280 ;
        RECT 521.370 0.155 525.130 4.280 ;
        RECT 525.970 0.155 529.730 4.280 ;
        RECT 530.570 0.155 534.330 4.280 ;
        RECT 535.170 0.155 538.010 4.280 ;
        RECT 538.850 0.155 542.610 4.280 ;
        RECT 543.450 0.155 547.210 4.280 ;
        RECT 548.050 0.155 551.810 4.280 ;
        RECT 552.650 0.155 555.490 4.280 ;
        RECT 556.330 0.155 560.090 4.280 ;
        RECT 560.930 0.155 564.690 4.280 ;
        RECT 565.530 0.155 569.290 4.280 ;
        RECT 570.130 0.155 572.970 4.280 ;
        RECT 573.810 0.155 577.570 4.280 ;
        RECT 578.410 0.155 582.170 4.280 ;
        RECT 583.010 0.155 586.770 4.280 ;
        RECT 587.610 0.155 590.450 4.280 ;
        RECT 591.290 0.155 595.050 4.280 ;
      LAYER met3 ;
        RECT 4.400 595.320 595.600 596.185 ;
        RECT 4.000 589.920 596.000 595.320 ;
        RECT 4.400 588.520 595.600 589.920 ;
        RECT 4.000 584.480 596.000 588.520 ;
        RECT 4.000 583.120 595.600 584.480 ;
        RECT 4.400 583.080 595.600 583.120 ;
        RECT 4.400 581.720 596.000 583.080 ;
        RECT 4.000 577.680 596.000 581.720 ;
        RECT 4.000 576.320 595.600 577.680 ;
        RECT 4.400 576.280 595.600 576.320 ;
        RECT 4.400 574.920 596.000 576.280 ;
        RECT 4.000 570.880 596.000 574.920 ;
        RECT 4.400 569.480 595.600 570.880 ;
        RECT 4.000 564.080 596.000 569.480 ;
        RECT 4.400 562.680 595.600 564.080 ;
        RECT 4.000 558.640 596.000 562.680 ;
        RECT 4.000 557.280 595.600 558.640 ;
        RECT 4.400 557.240 595.600 557.280 ;
        RECT 4.400 555.880 596.000 557.240 ;
        RECT 4.000 551.840 596.000 555.880 ;
        RECT 4.000 550.480 595.600 551.840 ;
        RECT 4.400 550.440 595.600 550.480 ;
        RECT 4.400 549.080 596.000 550.440 ;
        RECT 4.000 545.040 596.000 549.080 ;
        RECT 4.400 543.640 595.600 545.040 ;
        RECT 4.000 538.240 596.000 543.640 ;
        RECT 4.400 536.840 595.600 538.240 ;
        RECT 4.000 531.440 596.000 536.840 ;
        RECT 4.400 530.040 595.600 531.440 ;
        RECT 4.000 526.000 596.000 530.040 ;
        RECT 4.000 524.640 595.600 526.000 ;
        RECT 4.400 524.600 595.600 524.640 ;
        RECT 4.400 523.240 596.000 524.600 ;
        RECT 4.000 519.200 596.000 523.240 ;
        RECT 4.400 517.800 595.600 519.200 ;
        RECT 4.000 512.400 596.000 517.800 ;
        RECT 4.400 511.000 595.600 512.400 ;
        RECT 4.000 505.600 596.000 511.000 ;
        RECT 4.400 504.200 595.600 505.600 ;
        RECT 4.000 500.160 596.000 504.200 ;
        RECT 4.000 498.800 595.600 500.160 ;
        RECT 4.400 498.760 595.600 498.800 ;
        RECT 4.400 497.400 596.000 498.760 ;
        RECT 4.000 493.360 596.000 497.400 ;
        RECT 4.000 492.000 595.600 493.360 ;
        RECT 4.400 491.960 595.600 492.000 ;
        RECT 4.400 490.600 596.000 491.960 ;
        RECT 4.000 486.560 596.000 490.600 ;
        RECT 4.400 485.160 595.600 486.560 ;
        RECT 4.000 479.760 596.000 485.160 ;
        RECT 4.400 478.360 595.600 479.760 ;
        RECT 4.000 474.320 596.000 478.360 ;
        RECT 4.000 472.960 595.600 474.320 ;
        RECT 4.400 472.920 595.600 472.960 ;
        RECT 4.400 471.560 596.000 472.920 ;
        RECT 4.000 467.520 596.000 471.560 ;
        RECT 4.000 466.160 595.600 467.520 ;
        RECT 4.400 466.120 595.600 466.160 ;
        RECT 4.400 464.760 596.000 466.120 ;
        RECT 4.000 460.720 596.000 464.760 ;
        RECT 4.400 459.320 595.600 460.720 ;
        RECT 4.000 453.920 596.000 459.320 ;
        RECT 4.400 452.520 595.600 453.920 ;
        RECT 4.000 448.480 596.000 452.520 ;
        RECT 4.000 447.120 595.600 448.480 ;
        RECT 4.400 447.080 595.600 447.120 ;
        RECT 4.400 445.720 596.000 447.080 ;
        RECT 4.000 441.680 596.000 445.720 ;
        RECT 4.000 440.320 595.600 441.680 ;
        RECT 4.400 440.280 595.600 440.320 ;
        RECT 4.400 438.920 596.000 440.280 ;
        RECT 4.000 434.880 596.000 438.920 ;
        RECT 4.400 433.480 595.600 434.880 ;
        RECT 4.000 428.080 596.000 433.480 ;
        RECT 4.400 426.680 595.600 428.080 ;
        RECT 4.000 422.640 596.000 426.680 ;
        RECT 4.000 421.280 595.600 422.640 ;
        RECT 4.400 421.240 595.600 421.280 ;
        RECT 4.400 419.880 596.000 421.240 ;
        RECT 4.000 415.840 596.000 419.880 ;
        RECT 4.000 414.480 595.600 415.840 ;
        RECT 4.400 414.440 595.600 414.480 ;
        RECT 4.400 413.080 596.000 414.440 ;
        RECT 4.000 409.040 596.000 413.080 ;
        RECT 4.400 407.640 595.600 409.040 ;
        RECT 4.000 402.240 596.000 407.640 ;
        RECT 4.400 400.840 595.600 402.240 ;
        RECT 4.000 395.440 596.000 400.840 ;
        RECT 4.400 394.040 595.600 395.440 ;
        RECT 4.000 390.000 596.000 394.040 ;
        RECT 4.000 388.640 595.600 390.000 ;
        RECT 4.400 388.600 595.600 388.640 ;
        RECT 4.400 387.240 596.000 388.600 ;
        RECT 4.000 383.200 596.000 387.240 ;
        RECT 4.000 381.840 595.600 383.200 ;
        RECT 4.400 381.800 595.600 381.840 ;
        RECT 4.400 380.440 596.000 381.800 ;
        RECT 4.000 376.400 596.000 380.440 ;
        RECT 4.400 375.000 595.600 376.400 ;
        RECT 4.000 369.600 596.000 375.000 ;
        RECT 4.400 368.200 595.600 369.600 ;
        RECT 4.000 364.160 596.000 368.200 ;
        RECT 4.000 362.800 595.600 364.160 ;
        RECT 4.400 362.760 595.600 362.800 ;
        RECT 4.400 361.400 596.000 362.760 ;
        RECT 4.000 357.360 596.000 361.400 ;
        RECT 4.000 356.000 595.600 357.360 ;
        RECT 4.400 355.960 595.600 356.000 ;
        RECT 4.400 354.600 596.000 355.960 ;
        RECT 4.000 350.560 596.000 354.600 ;
        RECT 4.400 349.160 595.600 350.560 ;
        RECT 4.000 343.760 596.000 349.160 ;
        RECT 4.400 342.360 595.600 343.760 ;
        RECT 4.000 338.320 596.000 342.360 ;
        RECT 4.000 336.960 595.600 338.320 ;
        RECT 4.400 336.920 595.600 336.960 ;
        RECT 4.400 335.560 596.000 336.920 ;
        RECT 4.000 331.520 596.000 335.560 ;
        RECT 4.000 330.160 595.600 331.520 ;
        RECT 4.400 330.120 595.600 330.160 ;
        RECT 4.400 328.760 596.000 330.120 ;
        RECT 4.000 324.720 596.000 328.760 ;
        RECT 4.400 323.320 595.600 324.720 ;
        RECT 4.000 317.920 596.000 323.320 ;
        RECT 4.400 316.520 595.600 317.920 ;
        RECT 4.000 312.480 596.000 316.520 ;
        RECT 4.000 311.120 595.600 312.480 ;
        RECT 4.400 311.080 595.600 311.120 ;
        RECT 4.400 309.720 596.000 311.080 ;
        RECT 4.000 305.680 596.000 309.720 ;
        RECT 4.000 304.320 595.600 305.680 ;
        RECT 4.400 304.280 595.600 304.320 ;
        RECT 4.400 302.920 596.000 304.280 ;
        RECT 4.000 298.880 596.000 302.920 ;
        RECT 4.400 297.480 595.600 298.880 ;
        RECT 4.000 292.080 596.000 297.480 ;
        RECT 4.400 290.680 595.600 292.080 ;
        RECT 4.000 286.640 596.000 290.680 ;
        RECT 4.000 285.280 595.600 286.640 ;
        RECT 4.400 285.240 595.600 285.280 ;
        RECT 4.400 283.880 596.000 285.240 ;
        RECT 4.000 279.840 596.000 283.880 ;
        RECT 4.000 278.480 595.600 279.840 ;
        RECT 4.400 278.440 595.600 278.480 ;
        RECT 4.400 277.080 596.000 278.440 ;
        RECT 4.000 273.040 596.000 277.080 ;
        RECT 4.400 271.640 595.600 273.040 ;
        RECT 4.000 266.240 596.000 271.640 ;
        RECT 4.400 264.840 595.600 266.240 ;
        RECT 4.000 259.440 596.000 264.840 ;
        RECT 4.400 258.040 595.600 259.440 ;
        RECT 4.000 254.000 596.000 258.040 ;
        RECT 4.000 252.640 595.600 254.000 ;
        RECT 4.400 252.600 595.600 252.640 ;
        RECT 4.400 251.240 596.000 252.600 ;
        RECT 4.000 247.200 596.000 251.240 ;
        RECT 4.000 245.840 595.600 247.200 ;
        RECT 4.400 245.800 595.600 245.840 ;
        RECT 4.400 244.440 596.000 245.800 ;
        RECT 4.000 240.400 596.000 244.440 ;
        RECT 4.400 239.000 595.600 240.400 ;
        RECT 4.000 233.600 596.000 239.000 ;
        RECT 4.400 232.200 595.600 233.600 ;
        RECT 4.000 228.160 596.000 232.200 ;
        RECT 4.000 226.800 595.600 228.160 ;
        RECT 4.400 226.760 595.600 226.800 ;
        RECT 4.400 225.400 596.000 226.760 ;
        RECT 4.000 221.360 596.000 225.400 ;
        RECT 4.000 220.000 595.600 221.360 ;
        RECT 4.400 219.960 595.600 220.000 ;
        RECT 4.400 218.600 596.000 219.960 ;
        RECT 4.000 214.560 596.000 218.600 ;
        RECT 4.400 213.160 595.600 214.560 ;
        RECT 4.000 207.760 596.000 213.160 ;
        RECT 4.400 206.360 595.600 207.760 ;
        RECT 4.000 202.320 596.000 206.360 ;
        RECT 4.000 200.960 595.600 202.320 ;
        RECT 4.400 200.920 595.600 200.960 ;
        RECT 4.400 199.560 596.000 200.920 ;
        RECT 4.000 195.520 596.000 199.560 ;
        RECT 4.000 194.160 595.600 195.520 ;
        RECT 4.400 194.120 595.600 194.160 ;
        RECT 4.400 192.760 596.000 194.120 ;
        RECT 4.000 188.720 596.000 192.760 ;
        RECT 4.400 187.320 595.600 188.720 ;
        RECT 4.000 181.920 596.000 187.320 ;
        RECT 4.400 180.520 595.600 181.920 ;
        RECT 4.000 176.480 596.000 180.520 ;
        RECT 4.000 175.120 595.600 176.480 ;
        RECT 4.400 175.080 595.600 175.120 ;
        RECT 4.400 173.720 596.000 175.080 ;
        RECT 4.000 169.680 596.000 173.720 ;
        RECT 4.000 168.320 595.600 169.680 ;
        RECT 4.400 168.280 595.600 168.320 ;
        RECT 4.400 166.920 596.000 168.280 ;
        RECT 4.000 162.880 596.000 166.920 ;
        RECT 4.400 161.480 595.600 162.880 ;
        RECT 4.000 156.080 596.000 161.480 ;
        RECT 4.400 154.680 595.600 156.080 ;
        RECT 4.000 150.640 596.000 154.680 ;
        RECT 4.000 149.280 595.600 150.640 ;
        RECT 4.400 149.240 595.600 149.280 ;
        RECT 4.400 147.880 596.000 149.240 ;
        RECT 4.000 143.840 596.000 147.880 ;
        RECT 4.000 142.480 595.600 143.840 ;
        RECT 4.400 142.440 595.600 142.480 ;
        RECT 4.400 141.080 596.000 142.440 ;
        RECT 4.000 137.040 596.000 141.080 ;
        RECT 4.400 135.640 595.600 137.040 ;
        RECT 4.000 130.240 596.000 135.640 ;
        RECT 4.400 128.840 595.600 130.240 ;
        RECT 4.000 123.440 596.000 128.840 ;
        RECT 4.400 122.040 595.600 123.440 ;
        RECT 4.000 118.000 596.000 122.040 ;
        RECT 4.000 116.640 595.600 118.000 ;
        RECT 4.400 116.600 595.600 116.640 ;
        RECT 4.400 115.240 596.000 116.600 ;
        RECT 4.000 111.200 596.000 115.240 ;
        RECT 4.000 109.840 595.600 111.200 ;
        RECT 4.400 109.800 595.600 109.840 ;
        RECT 4.400 108.440 596.000 109.800 ;
        RECT 4.000 104.400 596.000 108.440 ;
        RECT 4.400 103.000 595.600 104.400 ;
        RECT 4.000 97.600 596.000 103.000 ;
        RECT 4.400 96.200 595.600 97.600 ;
        RECT 4.000 92.160 596.000 96.200 ;
        RECT 4.000 90.800 595.600 92.160 ;
        RECT 4.400 90.760 595.600 90.800 ;
        RECT 4.400 89.400 596.000 90.760 ;
        RECT 4.000 85.360 596.000 89.400 ;
        RECT 4.000 84.000 595.600 85.360 ;
        RECT 4.400 83.960 595.600 84.000 ;
        RECT 4.400 82.600 596.000 83.960 ;
        RECT 4.000 78.560 596.000 82.600 ;
        RECT 4.400 77.160 595.600 78.560 ;
        RECT 4.000 71.760 596.000 77.160 ;
        RECT 4.400 70.360 595.600 71.760 ;
        RECT 4.000 66.320 596.000 70.360 ;
        RECT 4.000 64.960 595.600 66.320 ;
        RECT 4.400 64.920 595.600 64.960 ;
        RECT 4.400 63.560 596.000 64.920 ;
        RECT 4.000 59.520 596.000 63.560 ;
        RECT 4.000 58.160 595.600 59.520 ;
        RECT 4.400 58.120 595.600 58.160 ;
        RECT 4.400 56.760 596.000 58.120 ;
        RECT 4.000 52.720 596.000 56.760 ;
        RECT 4.400 51.320 595.600 52.720 ;
        RECT 4.000 45.920 596.000 51.320 ;
        RECT 4.400 44.520 595.600 45.920 ;
        RECT 4.000 40.480 596.000 44.520 ;
        RECT 4.000 39.120 595.600 40.480 ;
        RECT 4.400 39.080 595.600 39.120 ;
        RECT 4.400 37.720 596.000 39.080 ;
        RECT 4.000 33.680 596.000 37.720 ;
        RECT 4.000 32.320 595.600 33.680 ;
        RECT 4.400 32.280 595.600 32.320 ;
        RECT 4.400 30.920 596.000 32.280 ;
        RECT 4.000 26.880 596.000 30.920 ;
        RECT 4.400 25.480 595.600 26.880 ;
        RECT 4.000 20.080 596.000 25.480 ;
        RECT 4.400 18.680 595.600 20.080 ;
        RECT 4.000 13.280 596.000 18.680 ;
        RECT 4.400 11.880 595.600 13.280 ;
        RECT 4.000 7.840 596.000 11.880 ;
        RECT 4.000 6.480 595.600 7.840 ;
        RECT 4.400 6.440 595.600 6.480 ;
        RECT 4.400 5.080 596.000 6.440 ;
        RECT 4.000 1.040 596.000 5.080 ;
        RECT 4.000 0.175 595.600 1.040 ;
      LAYER met4 ;
        RECT 189.815 38.935 251.040 435.025 ;
        RECT 253.440 38.935 327.840 435.025 ;
        RECT 330.240 38.935 404.505 435.025 ;
  END
END cache
END LIBRARY

