* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for chip_controller abstract view
.subckt chip_controller addr0_to_sram[0] addr0_to_sram[10] addr0_to_sram[11] addr0_to_sram[12]
+ addr0_to_sram[13] addr0_to_sram[14] addr0_to_sram[15] addr0_to_sram[16] addr0_to_sram[17]
+ addr0_to_sram[18] addr0_to_sram[19] addr0_to_sram[1] addr0_to_sram[2] addr0_to_sram[3]
+ addr0_to_sram[4] addr0_to_sram[5] addr0_to_sram[6] addr0_to_sram[7] addr0_to_sram[8]
+ addr0_to_sram[9] addr_in[0] addr_in[10] addr_in[11] addr_in[12] addr_in[13] addr_in[14]
+ addr_in[15] addr_in[16] addr_in[17] addr_in[18] addr_in[19] addr_in[1] addr_in[2]
+ addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in[8] addr_in[9] addr_to_core_mem[0]
+ addr_to_core_mem[10] addr_to_core_mem[11] addr_to_core_mem[12] addr_to_core_mem[13]
+ addr_to_core_mem[14] addr_to_core_mem[15] addr_to_core_mem[16] addr_to_core_mem[17]
+ addr_to_core_mem[18] addr_to_core_mem[19] addr_to_core_mem[1] addr_to_core_mem[2]
+ addr_to_core_mem[3] addr_to_core_mem[4] addr_to_core_mem[5] addr_to_core_mem[6]
+ addr_to_core_mem[7] addr_to_core_mem[8] addr_to_core_mem[9] clk core0_data_print[0]
+ core0_data_print[10] core0_data_print[11] core0_data_print[12] core0_data_print[13]
+ core0_data_print[14] core0_data_print[15] core0_data_print[16] core0_data_print[17]
+ core0_data_print[18] core0_data_print[19] core0_data_print[1] core0_data_print[20]
+ core0_data_print[21] core0_data_print[22] core0_data_print[23] core0_data_print[24]
+ core0_data_print[25] core0_data_print[26] core0_data_print[27] core0_data_print[28]
+ core0_data_print[29] core0_data_print[2] core0_data_print[30] core0_data_print[31]
+ core0_data_print[3] core0_data_print[4] core0_data_print[5] core0_data_print[6]
+ core0_data_print[7] core0_data_print[8] core0_data_print[9] csb0_to_sram data_out_to_core[0]
+ data_out_to_core[10] data_out_to_core[11] data_out_to_core[12] data_out_to_core[13]
+ data_out_to_core[14] data_out_to_core[15] data_out_to_core[16] data_out_to_core[17]
+ data_out_to_core[18] data_out_to_core[19] data_out_to_core[1] data_out_to_core[20]
+ data_out_to_core[21] data_out_to_core[22] data_out_to_core[23] data_out_to_core[24]
+ data_out_to_core[25] data_out_to_core[26] data_out_to_core[27] data_out_to_core[28]
+ data_out_to_core[29] data_out_to_core[2] data_out_to_core[30] data_out_to_core[31]
+ data_out_to_core[3] data_out_to_core[4] data_out_to_core[5] data_out_to_core[6]
+ data_out_to_core[7] data_out_to_core[8] data_out_to_core[9] data_to_core_mem[0]
+ data_to_core_mem[10] data_to_core_mem[11] data_to_core_mem[12] data_to_core_mem[13]
+ data_to_core_mem[14] data_to_core_mem[15] data_to_core_mem[16] data_to_core_mem[17]
+ data_to_core_mem[18] data_to_core_mem[19] data_to_core_mem[1] data_to_core_mem[20]
+ data_to_core_mem[21] data_to_core_mem[22] data_to_core_mem[23] data_to_core_mem[24]
+ data_to_core_mem[25] data_to_core_mem[26] data_to_core_mem[27] data_to_core_mem[28]
+ data_to_core_mem[29] data_to_core_mem[2] data_to_core_mem[30] data_to_core_mem[31]
+ data_to_core_mem[3] data_to_core_mem[4] data_to_core_mem[5] data_to_core_mem[6]
+ data_to_core_mem[7] data_to_core_mem[8] data_to_core_mem[9] din0_to_sram[0] din0_to_sram[10]
+ din0_to_sram[11] din0_to_sram[12] din0_to_sram[13] din0_to_sram[14] din0_to_sram[15]
+ din0_to_sram[16] din0_to_sram[17] din0_to_sram[18] din0_to_sram[19] din0_to_sram[1]
+ din0_to_sram[20] din0_to_sram[21] din0_to_sram[22] din0_to_sram[23] din0_to_sram[24]
+ din0_to_sram[25] din0_to_sram[26] din0_to_sram[27] din0_to_sram[28] din0_to_sram[29]
+ din0_to_sram[2] din0_to_sram[30] din0_to_sram[31] din0_to_sram[3] din0_to_sram[4]
+ din0_to_sram[5] din0_to_sram[6] din0_to_sram[7] din0_to_sram[8] din0_to_sram[9]
+ dout0_to_sram[0] dout0_to_sram[10] dout0_to_sram[11] dout0_to_sram[12] dout0_to_sram[13]
+ dout0_to_sram[14] dout0_to_sram[15] dout0_to_sram[16] dout0_to_sram[17] dout0_to_sram[18]
+ dout0_to_sram[19] dout0_to_sram[1] dout0_to_sram[20] dout0_to_sram[21] dout0_to_sram[22]
+ dout0_to_sram[23] dout0_to_sram[24] dout0_to_sram[25] dout0_to_sram[26] dout0_to_sram[27]
+ dout0_to_sram[28] dout0_to_sram[29] dout0_to_sram[2] dout0_to_sram[30] dout0_to_sram[31]
+ dout0_to_sram[3] dout0_to_sram[4] dout0_to_sram[5] dout0_to_sram[6] dout0_to_sram[7]
+ dout0_to_sram[8] dout0_to_sram[9] is_loading_memory_into_core is_ready_dataout_core0
+ is_ready_print_core0 la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] rd_data_out[0] rd_data_out[100] rd_data_out[101]
+ rd_data_out[102] rd_data_out[103] rd_data_out[104] rd_data_out[105] rd_data_out[106]
+ rd_data_out[107] rd_data_out[108] rd_data_out[109] rd_data_out[10] rd_data_out[110]
+ rd_data_out[111] rd_data_out[112] rd_data_out[113] rd_data_out[114] rd_data_out[115]
+ rd_data_out[116] rd_data_out[117] rd_data_out[118] rd_data_out[119] rd_data_out[11]
+ rd_data_out[120] rd_data_out[121] rd_data_out[122] rd_data_out[123] rd_data_out[124]
+ rd_data_out[125] rd_data_out[126] rd_data_out[127] rd_data_out[12] rd_data_out[13]
+ rd_data_out[14] rd_data_out[15] rd_data_out[16] rd_data_out[17] rd_data_out[18]
+ rd_data_out[19] rd_data_out[1] rd_data_out[20] rd_data_out[21] rd_data_out[22] rd_data_out[23]
+ rd_data_out[24] rd_data_out[25] rd_data_out[26] rd_data_out[27] rd_data_out[28]
+ rd_data_out[29] rd_data_out[2] rd_data_out[30] rd_data_out[31] rd_data_out[32] rd_data_out[33]
+ rd_data_out[34] rd_data_out[35] rd_data_out[36] rd_data_out[37] rd_data_out[38]
+ rd_data_out[39] rd_data_out[3] rd_data_out[40] rd_data_out[41] rd_data_out[42] rd_data_out[43]
+ rd_data_out[44] rd_data_out[45] rd_data_out[46] rd_data_out[47] rd_data_out[48]
+ rd_data_out[49] rd_data_out[4] rd_data_out[50] rd_data_out[51] rd_data_out[52] rd_data_out[53]
+ rd_data_out[54] rd_data_out[55] rd_data_out[56] rd_data_out[57] rd_data_out[58]
+ rd_data_out[59] rd_data_out[5] rd_data_out[60] rd_data_out[61] rd_data_out[62] rd_data_out[63]
+ rd_data_out[64] rd_data_out[65] rd_data_out[66] rd_data_out[67] rd_data_out[68]
+ rd_data_out[69] rd_data_out[6] rd_data_out[70] rd_data_out[71] rd_data_out[72] rd_data_out[73]
+ rd_data_out[74] rd_data_out[75] rd_data_out[76] rd_data_out[77] rd_data_out[78]
+ rd_data_out[79] rd_data_out[7] rd_data_out[80] rd_data_out[81] rd_data_out[82] rd_data_out[83]
+ rd_data_out[84] rd_data_out[85] rd_data_out[86] rd_data_out[87] rd_data_out[88]
+ rd_data_out[89] rd_data_out[8] rd_data_out[90] rd_data_out[91] rd_data_out[92] rd_data_out[93]
+ rd_data_out[94] rd_data_out[95] rd_data_out[96] rd_data_out[97] rd_data_out[98]
+ rd_data_out[99] rd_data_out[9] read_enable_to_Elpis read_interactive_req_core0 read_value_to_Elpis[0]
+ read_value_to_Elpis[10] read_value_to_Elpis[11] read_value_to_Elpis[12] read_value_to_Elpis[13]
+ read_value_to_Elpis[14] read_value_to_Elpis[15] read_value_to_Elpis[16] read_value_to_Elpis[17]
+ read_value_to_Elpis[18] read_value_to_Elpis[19] read_value_to_Elpis[1] read_value_to_Elpis[20]
+ read_value_to_Elpis[21] read_value_to_Elpis[22] read_value_to_Elpis[23] read_value_to_Elpis[24]
+ read_value_to_Elpis[25] read_value_to_Elpis[26] read_value_to_Elpis[27] read_value_to_Elpis[28]
+ read_value_to_Elpis[29] read_value_to_Elpis[2] read_value_to_Elpis[30] read_value_to_Elpis[31]
+ read_value_to_Elpis[3] read_value_to_Elpis[4] read_value_to_Elpis[5] read_value_to_Elpis[6]
+ read_value_to_Elpis[7] read_value_to_Elpis[8] read_value_to_Elpis[9] ready req_out_core0
+ requested reset_core reset_mem_req rst spare_wen0_to_sram vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] we we_to_sram wr_data[0] wr_data[100] wr_data[101] wr_data[102] wr_data[103]
+ wr_data[104] wr_data[105] wr_data[106] wr_data[107] wr_data[108] wr_data[109] wr_data[10]
+ wr_data[110] wr_data[111] wr_data[112] wr_data[113] wr_data[114] wr_data[115] wr_data[116]
+ wr_data[117] wr_data[118] wr_data[119] wr_data[11] wr_data[120] wr_data[121] wr_data[122]
+ wr_data[123] wr_data[124] wr_data[125] wr_data[126] wr_data[127] wr_data[12] wr_data[13]
+ wr_data[14] wr_data[15] wr_data[16] wr_data[17] wr_data[18] wr_data[19] wr_data[1]
+ wr_data[20] wr_data[21] wr_data[22] wr_data[23] wr_data[24] wr_data[25] wr_data[26]
+ wr_data[27] wr_data[28] wr_data[29] wr_data[2] wr_data[30] wr_data[31] wr_data[32]
+ wr_data[33] wr_data[34] wr_data[35] wr_data[36] wr_data[37] wr_data[38] wr_data[39]
+ wr_data[3] wr_data[40] wr_data[41] wr_data[42] wr_data[43] wr_data[44] wr_data[45]
+ wr_data[46] wr_data[47] wr_data[48] wr_data[49] wr_data[4] wr_data[50] wr_data[51]
+ wr_data[52] wr_data[53] wr_data[54] wr_data[55] wr_data[56] wr_data[57] wr_data[58]
+ wr_data[59] wr_data[5] wr_data[60] wr_data[61] wr_data[62] wr_data[63] wr_data[64]
+ wr_data[65] wr_data[66] wr_data[67] wr_data[68] wr_data[69] wr_data[6] wr_data[70]
+ wr_data[71] wr_data[72] wr_data[73] wr_data[74] wr_data[75] wr_data[76] wr_data[77]
+ wr_data[78] wr_data[79] wr_data[7] wr_data[80] wr_data[81] wr_data[82] wr_data[83]
+ wr_data[84] wr_data[85] wr_data[86] wr_data[87] wr_data[88] wr_data[89] wr_data[8]
+ wr_data[90] wr_data[91] wr_data[92] wr_data[93] wr_data[94] wr_data[95] wr_data[96]
+ wr_data[97] wr_data[98] wr_data[99] wr_data[9]
.ends

* Black-box entry subcircuit for core abstract view
.subckt core clk data_from_mem[0] data_from_mem[100] data_from_mem[101] data_from_mem[102]
+ data_from_mem[103] data_from_mem[104] data_from_mem[105] data_from_mem[106] data_from_mem[107]
+ data_from_mem[108] data_from_mem[109] data_from_mem[10] data_from_mem[110] data_from_mem[111]
+ data_from_mem[112] data_from_mem[113] data_from_mem[114] data_from_mem[115] data_from_mem[116]
+ data_from_mem[117] data_from_mem[118] data_from_mem[119] data_from_mem[11] data_from_mem[120]
+ data_from_mem[121] data_from_mem[122] data_from_mem[123] data_from_mem[124] data_from_mem[125]
+ data_from_mem[126] data_from_mem[127] data_from_mem[12] data_from_mem[13] data_from_mem[14]
+ data_from_mem[15] data_from_mem[16] data_from_mem[17] data_from_mem[18] data_from_mem[19]
+ data_from_mem[1] data_from_mem[20] data_from_mem[21] data_from_mem[22] data_from_mem[23]
+ data_from_mem[24] data_from_mem[25] data_from_mem[26] data_from_mem[27] data_from_mem[28]
+ data_from_mem[29] data_from_mem[2] data_from_mem[30] data_from_mem[31] data_from_mem[32]
+ data_from_mem[33] data_from_mem[34] data_from_mem[35] data_from_mem[36] data_from_mem[37]
+ data_from_mem[38] data_from_mem[39] data_from_mem[3] data_from_mem[40] data_from_mem[41]
+ data_from_mem[42] data_from_mem[43] data_from_mem[44] data_from_mem[45] data_from_mem[46]
+ data_from_mem[47] data_from_mem[48] data_from_mem[49] data_from_mem[4] data_from_mem[50]
+ data_from_mem[51] data_from_mem[52] data_from_mem[53] data_from_mem[54] data_from_mem[55]
+ data_from_mem[56] data_from_mem[57] data_from_mem[58] data_from_mem[59] data_from_mem[5]
+ data_from_mem[60] data_from_mem[61] data_from_mem[62] data_from_mem[63] data_from_mem[64]
+ data_from_mem[65] data_from_mem[66] data_from_mem[67] data_from_mem[68] data_from_mem[69]
+ data_from_mem[6] data_from_mem[70] data_from_mem[71] data_from_mem[72] data_from_mem[73]
+ data_from_mem[74] data_from_mem[75] data_from_mem[76] data_from_mem[77] data_from_mem[78]
+ data_from_mem[79] data_from_mem[7] data_from_mem[80] data_from_mem[81] data_from_mem[82]
+ data_from_mem[83] data_from_mem[84] data_from_mem[85] data_from_mem[86] data_from_mem[87]
+ data_from_mem[88] data_from_mem[89] data_from_mem[8] data_from_mem[90] data_from_mem[91]
+ data_from_mem[92] data_from_mem[93] data_from_mem[94] data_from_mem[95] data_from_mem[96]
+ data_from_mem[97] data_from_mem[98] data_from_mem[99] data_from_mem[9] hex_out[0]
+ hex_out[10] hex_out[11] hex_out[12] hex_out[13] hex_out[14] hex_out[15] hex_out[16]
+ hex_out[17] hex_out[18] hex_out[19] hex_out[1] hex_out[20] hex_out[21] hex_out[22]
+ hex_out[23] hex_out[24] hex_out[25] hex_out[26] hex_out[27] hex_out[28] hex_out[29]
+ hex_out[2] hex_out[30] hex_out[31] hex_out[3] hex_out[4] hex_out[5] hex_out[6] hex_out[7]
+ hex_out[8] hex_out[9] hex_req is_mem_ready is_mem_req is_mem_req_reset is_memory_we
+ is_print_done mem_addr_out[0] mem_addr_out[10] mem_addr_out[11] mem_addr_out[12]
+ mem_addr_out[13] mem_addr_out[14] mem_addr_out[15] mem_addr_out[16] mem_addr_out[17]
+ mem_addr_out[18] mem_addr_out[19] mem_addr_out[1] mem_addr_out[2] mem_addr_out[3]
+ mem_addr_out[4] mem_addr_out[5] mem_addr_out[6] mem_addr_out[7] mem_addr_out[8]
+ mem_addr_out[9] mem_data_out[0] mem_data_out[100] mem_data_out[101] mem_data_out[102]
+ mem_data_out[103] mem_data_out[104] mem_data_out[105] mem_data_out[106] mem_data_out[107]
+ mem_data_out[108] mem_data_out[109] mem_data_out[10] mem_data_out[110] mem_data_out[111]
+ mem_data_out[112] mem_data_out[113] mem_data_out[114] mem_data_out[115] mem_data_out[116]
+ mem_data_out[117] mem_data_out[118] mem_data_out[119] mem_data_out[11] mem_data_out[120]
+ mem_data_out[121] mem_data_out[122] mem_data_out[123] mem_data_out[124] mem_data_out[125]
+ mem_data_out[126] mem_data_out[127] mem_data_out[12] mem_data_out[13] mem_data_out[14]
+ mem_data_out[15] mem_data_out[16] mem_data_out[17] mem_data_out[18] mem_data_out[19]
+ mem_data_out[1] mem_data_out[20] mem_data_out[21] mem_data_out[22] mem_data_out[23]
+ mem_data_out[24] mem_data_out[25] mem_data_out[26] mem_data_out[27] mem_data_out[28]
+ mem_data_out[29] mem_data_out[2] mem_data_out[30] mem_data_out[31] mem_data_out[32]
+ mem_data_out[33] mem_data_out[34] mem_data_out[35] mem_data_out[36] mem_data_out[37]
+ mem_data_out[38] mem_data_out[39] mem_data_out[3] mem_data_out[40] mem_data_out[41]
+ mem_data_out[42] mem_data_out[43] mem_data_out[44] mem_data_out[45] mem_data_out[46]
+ mem_data_out[47] mem_data_out[48] mem_data_out[49] mem_data_out[4] mem_data_out[50]
+ mem_data_out[51] mem_data_out[52] mem_data_out[53] mem_data_out[54] mem_data_out[55]
+ mem_data_out[56] mem_data_out[57] mem_data_out[58] mem_data_out[59] mem_data_out[5]
+ mem_data_out[60] mem_data_out[61] mem_data_out[62] mem_data_out[63] mem_data_out[64]
+ mem_data_out[65] mem_data_out[66] mem_data_out[67] mem_data_out[68] mem_data_out[69]
+ mem_data_out[6] mem_data_out[70] mem_data_out[71] mem_data_out[72] mem_data_out[73]
+ mem_data_out[74] mem_data_out[75] mem_data_out[76] mem_data_out[77] mem_data_out[78]
+ mem_data_out[79] mem_data_out[7] mem_data_out[80] mem_data_out[81] mem_data_out[82]
+ mem_data_out[83] mem_data_out[84] mem_data_out[85] mem_data_out[86] mem_data_out[87]
+ mem_data_out[88] mem_data_out[89] mem_data_out[8] mem_data_out[90] mem_data_out[91]
+ mem_data_out[92] mem_data_out[93] mem_data_out[94] mem_data_out[95] mem_data_out[96]
+ mem_data_out[97] mem_data_out[98] mem_data_out[99] mem_data_out[9] read_interactive_ready
+ read_interactive_req read_interactive_value[0] read_interactive_value[10] read_interactive_value[11]
+ read_interactive_value[12] read_interactive_value[13] read_interactive_value[14]
+ read_interactive_value[15] read_interactive_value[16] read_interactive_value[17]
+ read_interactive_value[18] read_interactive_value[19] read_interactive_value[1]
+ read_interactive_value[20] read_interactive_value[21] read_interactive_value[22]
+ read_interactive_value[23] read_interactive_value[24] read_interactive_value[25]
+ read_interactive_value[26] read_interactive_value[27] read_interactive_value[28]
+ read_interactive_value[29] read_interactive_value[2] read_interactive_value[30]
+ read_interactive_value[31] read_interactive_value[3] read_interactive_value[4] read_interactive_value[5]
+ read_interactive_value[6] read_interactive_value[7] read_interactive_value[8] read_interactive_value[9]
+ rst vccd1 vssd1
.ends

* Black-box entry subcircuit for custom_sram abstract view
.subckt custom_sram a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16] a[17] a[18] a[19]
+ a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] a[9] clk csb0_to_sram d[0] d[10] d[11] d[12]
+ d[13] d[14] d[15] d[16] d[17] d[18] d[19] d[1] d[20] d[21] d[22] d[23] d[24] d[25]
+ d[26] d[27] d[28] d[29] d[2] d[30] d[31] d[3] d[4] d[5] d[6] d[7] d[8] d[9] q[0]
+ q[10] q[11] q[12] q[13] q[14] q[15] q[16] q[17] q[18] q[19] q[1] q[20] q[21] q[22]
+ q[23] q[24] q[25] q[26] q[27] q[28] q[29] q[2] q[30] q[31] q[3] q[4] q[5] q[6] q[7]
+ q[8] q[9] spare_wen0_to_sram vccd1 vssd1 we
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xchip_controller custom_sram/a[0] custom_sram/a[10] custom_sram/a[11] custom_sram/a[12]
+ custom_sram/a[13] custom_sram/a[14] custom_sram/a[15] custom_sram/a[16] custom_sram/a[17]
+ custom_sram/a[18] custom_sram/a[19] custom_sram/a[1] custom_sram/a[2] custom_sram/a[3]
+ custom_sram/a[4] custom_sram/a[5] custom_sram/a[6] custom_sram/a[7] custom_sram/a[8]
+ custom_sram/a[9] core0/mem_addr_out[0] core0/mem_addr_out[10] core0/mem_addr_out[11]
+ core0/mem_addr_out[12] core0/mem_addr_out[13] core0/mem_addr_out[14] core0/mem_addr_out[15]
+ core0/mem_addr_out[16] core0/mem_addr_out[17] core0/mem_addr_out[18] core0/mem_addr_out[19]
+ core0/mem_addr_out[1] core0/mem_addr_out[2] core0/mem_addr_out[3] core0/mem_addr_out[4]
+ core0/mem_addr_out[5] core0/mem_addr_out[6] core0/mem_addr_out[7] core0/mem_addr_out[8]
+ core0/mem_addr_out[9] chip_controller/addr_to_core_mem[0] chip_controller/addr_to_core_mem[10]
+ chip_controller/addr_to_core_mem[11] chip_controller/addr_to_core_mem[12] chip_controller/addr_to_core_mem[13]
+ chip_controller/addr_to_core_mem[14] chip_controller/addr_to_core_mem[15] chip_controller/addr_to_core_mem[16]
+ chip_controller/addr_to_core_mem[17] chip_controller/addr_to_core_mem[18] chip_controller/addr_to_core_mem[19]
+ chip_controller/addr_to_core_mem[1] chip_controller/addr_to_core_mem[2] chip_controller/addr_to_core_mem[3]
+ chip_controller/addr_to_core_mem[4] chip_controller/addr_to_core_mem[5] chip_controller/addr_to_core_mem[6]
+ chip_controller/addr_to_core_mem[7] chip_controller/addr_to_core_mem[8] chip_controller/addr_to_core_mem[9]
+ core0/clk core0/hex_out[0] core0/hex_out[10] core0/hex_out[11] core0/hex_out[12]
+ core0/hex_out[13] core0/hex_out[14] core0/hex_out[15] core0/hex_out[16] core0/hex_out[17]
+ core0/hex_out[18] core0/hex_out[19] core0/hex_out[1] core0/hex_out[20] core0/hex_out[21]
+ core0/hex_out[22] core0/hex_out[23] core0/hex_out[24] core0/hex_out[25] core0/hex_out[26]
+ core0/hex_out[27] core0/hex_out[28] core0/hex_out[29] core0/hex_out[2] core0/hex_out[30]
+ core0/hex_out[31] core0/hex_out[3] core0/hex_out[4] core0/hex_out[5] core0/hex_out[6]
+ core0/hex_out[7] core0/hex_out[8] core0/hex_out[9] custom_sram/csb0_to_sram core0/read_interactive_value[0]
+ core0/read_interactive_value[10] core0/read_interactive_value[11] core0/read_interactive_value[12]
+ core0/read_interactive_value[13] core0/read_interactive_value[14] core0/read_interactive_value[15]
+ core0/read_interactive_value[16] core0/read_interactive_value[17] core0/read_interactive_value[18]
+ core0/read_interactive_value[19] core0/read_interactive_value[1] core0/read_interactive_value[20]
+ core0/read_interactive_value[21] core0/read_interactive_value[22] core0/read_interactive_value[23]
+ core0/read_interactive_value[24] core0/read_interactive_value[25] core0/read_interactive_value[26]
+ core0/read_interactive_value[27] core0/read_interactive_value[28] core0/read_interactive_value[29]
+ core0/read_interactive_value[2] core0/read_interactive_value[30] core0/read_interactive_value[31]
+ core0/read_interactive_value[3] core0/read_interactive_value[4] core0/read_interactive_value[5]
+ core0/read_interactive_value[6] core0/read_interactive_value[7] core0/read_interactive_value[8]
+ core0/read_interactive_value[9] chip_controller/data_to_core_mem[0] chip_controller/data_to_core_mem[10]
+ chip_controller/data_to_core_mem[11] chip_controller/data_to_core_mem[12] chip_controller/data_to_core_mem[13]
+ chip_controller/data_to_core_mem[14] chip_controller/data_to_core_mem[15] chip_controller/data_to_core_mem[16]
+ chip_controller/data_to_core_mem[17] chip_controller/data_to_core_mem[18] chip_controller/data_to_core_mem[19]
+ chip_controller/data_to_core_mem[1] chip_controller/data_to_core_mem[20] chip_controller/data_to_core_mem[21]
+ chip_controller/data_to_core_mem[22] chip_controller/data_to_core_mem[23] chip_controller/data_to_core_mem[24]
+ chip_controller/data_to_core_mem[25] chip_controller/data_to_core_mem[26] chip_controller/data_to_core_mem[27]
+ chip_controller/data_to_core_mem[28] chip_controller/data_to_core_mem[29] chip_controller/data_to_core_mem[2]
+ chip_controller/data_to_core_mem[30] chip_controller/data_to_core_mem[31] chip_controller/data_to_core_mem[3]
+ chip_controller/data_to_core_mem[4] chip_controller/data_to_core_mem[5] chip_controller/data_to_core_mem[6]
+ chip_controller/data_to_core_mem[7] chip_controller/data_to_core_mem[8] chip_controller/data_to_core_mem[9]
+ custom_sram/d[0] custom_sram/d[10] custom_sram/d[11] custom_sram/d[12] custom_sram/d[13]
+ custom_sram/d[14] custom_sram/d[15] custom_sram/d[16] custom_sram/d[17] custom_sram/d[18]
+ custom_sram/d[19] custom_sram/d[1] custom_sram/d[20] custom_sram/d[21] custom_sram/d[22]
+ custom_sram/d[23] custom_sram/d[24] custom_sram/d[25] custom_sram/d[26] custom_sram/d[27]
+ custom_sram/d[28] custom_sram/d[29] custom_sram/d[2] custom_sram/d[30] custom_sram/d[31]
+ custom_sram/d[3] custom_sram/d[4] custom_sram/d[5] custom_sram/d[6] custom_sram/d[7]
+ custom_sram/d[8] custom_sram/d[9] custom_sram/q[0] custom_sram/q[10] custom_sram/q[11]
+ custom_sram/q[12] custom_sram/q[13] custom_sram/q[14] custom_sram/q[15] custom_sram/q[16]
+ custom_sram/q[17] custom_sram/q[18] custom_sram/q[19] custom_sram/q[1] custom_sram/q[20]
+ custom_sram/q[21] custom_sram/q[22] custom_sram/q[23] custom_sram/q[24] custom_sram/q[25]
+ custom_sram/q[26] custom_sram/q[27] custom_sram/q[28] custom_sram/q[29] custom_sram/q[2]
+ custom_sram/q[30] custom_sram/q[31] custom_sram/q[3] custom_sram/q[4] custom_sram/q[5]
+ custom_sram/q[6] custom_sram/q[7] custom_sram/q[8] custom_sram/q[9] chip_controller/is_loading_memory_into_core
+ core0/read_interactive_ready core0/is_print_done la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] core0/data_from_mem[0] core0/data_from_mem[100]
+ core0/data_from_mem[101] core0/data_from_mem[102] core0/data_from_mem[103] core0/data_from_mem[104]
+ core0/data_from_mem[105] core0/data_from_mem[106] core0/data_from_mem[107] core0/data_from_mem[108]
+ core0/data_from_mem[109] core0/data_from_mem[10] core0/data_from_mem[110] core0/data_from_mem[111]
+ core0/data_from_mem[112] core0/data_from_mem[113] core0/data_from_mem[114] core0/data_from_mem[115]
+ core0/data_from_mem[116] core0/data_from_mem[117] core0/data_from_mem[118] core0/data_from_mem[119]
+ core0/data_from_mem[11] core0/data_from_mem[120] core0/data_from_mem[121] core0/data_from_mem[122]
+ core0/data_from_mem[123] core0/data_from_mem[124] core0/data_from_mem[125] core0/data_from_mem[126]
+ core0/data_from_mem[127] core0/data_from_mem[12] core0/data_from_mem[13] core0/data_from_mem[14]
+ core0/data_from_mem[15] core0/data_from_mem[16] core0/data_from_mem[17] core0/data_from_mem[18]
+ core0/data_from_mem[19] core0/data_from_mem[1] core0/data_from_mem[20] core0/data_from_mem[21]
+ core0/data_from_mem[22] core0/data_from_mem[23] core0/data_from_mem[24] core0/data_from_mem[25]
+ core0/data_from_mem[26] core0/data_from_mem[27] core0/data_from_mem[28] core0/data_from_mem[29]
+ core0/data_from_mem[2] core0/data_from_mem[30] core0/data_from_mem[31] core0/data_from_mem[32]
+ core0/data_from_mem[33] core0/data_from_mem[34] core0/data_from_mem[35] core0/data_from_mem[36]
+ core0/data_from_mem[37] core0/data_from_mem[38] core0/data_from_mem[39] core0/data_from_mem[3]
+ core0/data_from_mem[40] core0/data_from_mem[41] core0/data_from_mem[42] core0/data_from_mem[43]
+ core0/data_from_mem[44] core0/data_from_mem[45] core0/data_from_mem[46] core0/data_from_mem[47]
+ core0/data_from_mem[48] core0/data_from_mem[49] core0/data_from_mem[4] core0/data_from_mem[50]
+ core0/data_from_mem[51] core0/data_from_mem[52] core0/data_from_mem[53] core0/data_from_mem[54]
+ core0/data_from_mem[55] core0/data_from_mem[56] core0/data_from_mem[57] core0/data_from_mem[58]
+ core0/data_from_mem[59] core0/data_from_mem[5] core0/data_from_mem[60] core0/data_from_mem[61]
+ core0/data_from_mem[62] core0/data_from_mem[63] core0/data_from_mem[64] core0/data_from_mem[65]
+ core0/data_from_mem[66] core0/data_from_mem[67] core0/data_from_mem[68] core0/data_from_mem[69]
+ core0/data_from_mem[6] core0/data_from_mem[70] core0/data_from_mem[71] core0/data_from_mem[72]
+ core0/data_from_mem[73] core0/data_from_mem[74] core0/data_from_mem[75] core0/data_from_mem[76]
+ core0/data_from_mem[77] core0/data_from_mem[78] core0/data_from_mem[79] core0/data_from_mem[7]
+ core0/data_from_mem[80] core0/data_from_mem[81] core0/data_from_mem[82] core0/data_from_mem[83]
+ core0/data_from_mem[84] core0/data_from_mem[85] core0/data_from_mem[86] core0/data_from_mem[87]
+ core0/data_from_mem[88] core0/data_from_mem[89] core0/data_from_mem[8] core0/data_from_mem[90]
+ core0/data_from_mem[91] core0/data_from_mem[92] core0/data_from_mem[93] core0/data_from_mem[94]
+ core0/data_from_mem[95] core0/data_from_mem[96] core0/data_from_mem[97] core0/data_from_mem[98]
+ core0/data_from_mem[99] core0/data_from_mem[9] chip_controller/read_enable_to_Elpis
+ core0/read_interactive_req chip_controller/read_value_to_Elpis[0] chip_controller/read_value_to_Elpis[10]
+ chip_controller/read_value_to_Elpis[11] chip_controller/read_value_to_Elpis[12]
+ chip_controller/read_value_to_Elpis[13] chip_controller/read_value_to_Elpis[14]
+ chip_controller/read_value_to_Elpis[15] chip_controller/read_value_to_Elpis[16]
+ chip_controller/read_value_to_Elpis[17] chip_controller/read_value_to_Elpis[18]
+ chip_controller/read_value_to_Elpis[19] chip_controller/read_value_to_Elpis[1] chip_controller/read_value_to_Elpis[20]
+ chip_controller/read_value_to_Elpis[21] chip_controller/read_value_to_Elpis[22]
+ chip_controller/read_value_to_Elpis[23] chip_controller/read_value_to_Elpis[24]
+ chip_controller/read_value_to_Elpis[25] chip_controller/read_value_to_Elpis[26]
+ chip_controller/read_value_to_Elpis[27] chip_controller/read_value_to_Elpis[28]
+ chip_controller/read_value_to_Elpis[29] chip_controller/read_value_to_Elpis[2] chip_controller/read_value_to_Elpis[30]
+ chip_controller/read_value_to_Elpis[31] chip_controller/read_value_to_Elpis[3] chip_controller/read_value_to_Elpis[4]
+ chip_controller/read_value_to_Elpis[5] chip_controller/read_value_to_Elpis[6] chip_controller/read_value_to_Elpis[7]
+ chip_controller/read_value_to_Elpis[8] chip_controller/read_value_to_Elpis[9] core0/is_mem_ready
+ core0/hex_req core0/is_mem_req core0/rst core0/is_mem_req_reset chip_controller/rst
+ custom_sram/spare_wen0_to_sram vccd1 vssd1 wb_clk_i wb_rst_i wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] core0/is_memory_we
+ custom_sram/we core0/mem_data_out[0] core0/mem_data_out[100] core0/mem_data_out[101]
+ core0/mem_data_out[102] core0/mem_data_out[103] core0/mem_data_out[104] core0/mem_data_out[105]
+ core0/mem_data_out[106] core0/mem_data_out[107] core0/mem_data_out[108] core0/mem_data_out[109]
+ core0/mem_data_out[10] core0/mem_data_out[110] core0/mem_data_out[111] core0/mem_data_out[112]
+ core0/mem_data_out[113] core0/mem_data_out[114] core0/mem_data_out[115] core0/mem_data_out[116]
+ core0/mem_data_out[117] core0/mem_data_out[118] core0/mem_data_out[119] core0/mem_data_out[11]
+ core0/mem_data_out[120] core0/mem_data_out[121] core0/mem_data_out[122] core0/mem_data_out[123]
+ core0/mem_data_out[124] core0/mem_data_out[125] core0/mem_data_out[126] core0/mem_data_out[127]
+ core0/mem_data_out[12] core0/mem_data_out[13] core0/mem_data_out[14] core0/mem_data_out[15]
+ core0/mem_data_out[16] core0/mem_data_out[17] core0/mem_data_out[18] core0/mem_data_out[19]
+ core0/mem_data_out[1] core0/mem_data_out[20] core0/mem_data_out[21] core0/mem_data_out[22]
+ core0/mem_data_out[23] core0/mem_data_out[24] core0/mem_data_out[25] core0/mem_data_out[26]
+ core0/mem_data_out[27] core0/mem_data_out[28] core0/mem_data_out[29] core0/mem_data_out[2]
+ core0/mem_data_out[30] core0/mem_data_out[31] core0/mem_data_out[32] core0/mem_data_out[33]
+ core0/mem_data_out[34] core0/mem_data_out[35] core0/mem_data_out[36] core0/mem_data_out[37]
+ core0/mem_data_out[38] core0/mem_data_out[39] core0/mem_data_out[3] core0/mem_data_out[40]
+ core0/mem_data_out[41] core0/mem_data_out[42] core0/mem_data_out[43] core0/mem_data_out[44]
+ core0/mem_data_out[45] core0/mem_data_out[46] core0/mem_data_out[47] core0/mem_data_out[48]
+ core0/mem_data_out[49] core0/mem_data_out[4] core0/mem_data_out[50] core0/mem_data_out[51]
+ core0/mem_data_out[52] core0/mem_data_out[53] core0/mem_data_out[54] core0/mem_data_out[55]
+ core0/mem_data_out[56] core0/mem_data_out[57] core0/mem_data_out[58] core0/mem_data_out[59]
+ core0/mem_data_out[5] core0/mem_data_out[60] core0/mem_data_out[61] core0/mem_data_out[62]
+ core0/mem_data_out[63] core0/mem_data_out[64] core0/mem_data_out[65] core0/mem_data_out[66]
+ core0/mem_data_out[67] core0/mem_data_out[68] core0/mem_data_out[69] core0/mem_data_out[6]
+ core0/mem_data_out[70] core0/mem_data_out[71] core0/mem_data_out[72] core0/mem_data_out[73]
+ core0/mem_data_out[74] core0/mem_data_out[75] core0/mem_data_out[76] core0/mem_data_out[77]
+ core0/mem_data_out[78] core0/mem_data_out[79] core0/mem_data_out[7] core0/mem_data_out[80]
+ core0/mem_data_out[81] core0/mem_data_out[82] core0/mem_data_out[83] core0/mem_data_out[84]
+ core0/mem_data_out[85] core0/mem_data_out[86] core0/mem_data_out[87] core0/mem_data_out[88]
+ core0/mem_data_out[89] core0/mem_data_out[8] core0/mem_data_out[90] core0/mem_data_out[91]
+ core0/mem_data_out[92] core0/mem_data_out[93] core0/mem_data_out[94] core0/mem_data_out[95]
+ core0/mem_data_out[96] core0/mem_data_out[97] core0/mem_data_out[98] core0/mem_data_out[99]
+ core0/mem_data_out[9] chip_controller
Xcore0 core0/clk core0/data_from_mem[0] core0/data_from_mem[100] core0/data_from_mem[101]
+ core0/data_from_mem[102] core0/data_from_mem[103] core0/data_from_mem[104] core0/data_from_mem[105]
+ core0/data_from_mem[106] core0/data_from_mem[107] core0/data_from_mem[108] core0/data_from_mem[109]
+ core0/data_from_mem[10] core0/data_from_mem[110] core0/data_from_mem[111] core0/data_from_mem[112]
+ core0/data_from_mem[113] core0/data_from_mem[114] core0/data_from_mem[115] core0/data_from_mem[116]
+ core0/data_from_mem[117] core0/data_from_mem[118] core0/data_from_mem[119] core0/data_from_mem[11]
+ core0/data_from_mem[120] core0/data_from_mem[121] core0/data_from_mem[122] core0/data_from_mem[123]
+ core0/data_from_mem[124] core0/data_from_mem[125] core0/data_from_mem[126] core0/data_from_mem[127]
+ core0/data_from_mem[12] core0/data_from_mem[13] core0/data_from_mem[14] core0/data_from_mem[15]
+ core0/data_from_mem[16] core0/data_from_mem[17] core0/data_from_mem[18] core0/data_from_mem[19]
+ core0/data_from_mem[1] core0/data_from_mem[20] core0/data_from_mem[21] core0/data_from_mem[22]
+ core0/data_from_mem[23] core0/data_from_mem[24] core0/data_from_mem[25] core0/data_from_mem[26]
+ core0/data_from_mem[27] core0/data_from_mem[28] core0/data_from_mem[29] core0/data_from_mem[2]
+ core0/data_from_mem[30] core0/data_from_mem[31] core0/data_from_mem[32] core0/data_from_mem[33]
+ core0/data_from_mem[34] core0/data_from_mem[35] core0/data_from_mem[36] core0/data_from_mem[37]
+ core0/data_from_mem[38] core0/data_from_mem[39] core0/data_from_mem[3] core0/data_from_mem[40]
+ core0/data_from_mem[41] core0/data_from_mem[42] core0/data_from_mem[43] core0/data_from_mem[44]
+ core0/data_from_mem[45] core0/data_from_mem[46] core0/data_from_mem[47] core0/data_from_mem[48]
+ core0/data_from_mem[49] core0/data_from_mem[4] core0/data_from_mem[50] core0/data_from_mem[51]
+ core0/data_from_mem[52] core0/data_from_mem[53] core0/data_from_mem[54] core0/data_from_mem[55]
+ core0/data_from_mem[56] core0/data_from_mem[57] core0/data_from_mem[58] core0/data_from_mem[59]
+ core0/data_from_mem[5] core0/data_from_mem[60] core0/data_from_mem[61] core0/data_from_mem[62]
+ core0/data_from_mem[63] core0/data_from_mem[64] core0/data_from_mem[65] core0/data_from_mem[66]
+ core0/data_from_mem[67] core0/data_from_mem[68] core0/data_from_mem[69] core0/data_from_mem[6]
+ core0/data_from_mem[70] core0/data_from_mem[71] core0/data_from_mem[72] core0/data_from_mem[73]
+ core0/data_from_mem[74] core0/data_from_mem[75] core0/data_from_mem[76] core0/data_from_mem[77]
+ core0/data_from_mem[78] core0/data_from_mem[79] core0/data_from_mem[7] core0/data_from_mem[80]
+ core0/data_from_mem[81] core0/data_from_mem[82] core0/data_from_mem[83] core0/data_from_mem[84]
+ core0/data_from_mem[85] core0/data_from_mem[86] core0/data_from_mem[87] core0/data_from_mem[88]
+ core0/data_from_mem[89] core0/data_from_mem[8] core0/data_from_mem[90] core0/data_from_mem[91]
+ core0/data_from_mem[92] core0/data_from_mem[93] core0/data_from_mem[94] core0/data_from_mem[95]
+ core0/data_from_mem[96] core0/data_from_mem[97] core0/data_from_mem[98] core0/data_from_mem[99]
+ core0/data_from_mem[9] core0/hex_out[0] core0/hex_out[10] core0/hex_out[11] core0/hex_out[12]
+ core0/hex_out[13] core0/hex_out[14] core0/hex_out[15] core0/hex_out[16] core0/hex_out[17]
+ core0/hex_out[18] core0/hex_out[19] core0/hex_out[1] core0/hex_out[20] core0/hex_out[21]
+ core0/hex_out[22] core0/hex_out[23] core0/hex_out[24] core0/hex_out[25] core0/hex_out[26]
+ core0/hex_out[27] core0/hex_out[28] core0/hex_out[29] core0/hex_out[2] core0/hex_out[30]
+ core0/hex_out[31] core0/hex_out[3] core0/hex_out[4] core0/hex_out[5] core0/hex_out[6]
+ core0/hex_out[7] core0/hex_out[8] core0/hex_out[9] core0/hex_req core0/is_mem_ready
+ core0/is_mem_req core0/is_mem_req_reset core0/is_memory_we core0/is_print_done core0/mem_addr_out[0]
+ core0/mem_addr_out[10] core0/mem_addr_out[11] core0/mem_addr_out[12] core0/mem_addr_out[13]
+ core0/mem_addr_out[14] core0/mem_addr_out[15] core0/mem_addr_out[16] core0/mem_addr_out[17]
+ core0/mem_addr_out[18] core0/mem_addr_out[19] core0/mem_addr_out[1] core0/mem_addr_out[2]
+ core0/mem_addr_out[3] core0/mem_addr_out[4] core0/mem_addr_out[5] core0/mem_addr_out[6]
+ core0/mem_addr_out[7] core0/mem_addr_out[8] core0/mem_addr_out[9] core0/mem_data_out[0]
+ core0/mem_data_out[100] core0/mem_data_out[101] core0/mem_data_out[102] core0/mem_data_out[103]
+ core0/mem_data_out[104] core0/mem_data_out[105] core0/mem_data_out[106] core0/mem_data_out[107]
+ core0/mem_data_out[108] core0/mem_data_out[109] core0/mem_data_out[10] core0/mem_data_out[110]
+ core0/mem_data_out[111] core0/mem_data_out[112] core0/mem_data_out[113] core0/mem_data_out[114]
+ core0/mem_data_out[115] core0/mem_data_out[116] core0/mem_data_out[117] core0/mem_data_out[118]
+ core0/mem_data_out[119] core0/mem_data_out[11] core0/mem_data_out[120] core0/mem_data_out[121]
+ core0/mem_data_out[122] core0/mem_data_out[123] core0/mem_data_out[124] core0/mem_data_out[125]
+ core0/mem_data_out[126] core0/mem_data_out[127] core0/mem_data_out[12] core0/mem_data_out[13]
+ core0/mem_data_out[14] core0/mem_data_out[15] core0/mem_data_out[16] core0/mem_data_out[17]
+ core0/mem_data_out[18] core0/mem_data_out[19] core0/mem_data_out[1] core0/mem_data_out[20]
+ core0/mem_data_out[21] core0/mem_data_out[22] core0/mem_data_out[23] core0/mem_data_out[24]
+ core0/mem_data_out[25] core0/mem_data_out[26] core0/mem_data_out[27] core0/mem_data_out[28]
+ core0/mem_data_out[29] core0/mem_data_out[2] core0/mem_data_out[30] core0/mem_data_out[31]
+ core0/mem_data_out[32] core0/mem_data_out[33] core0/mem_data_out[34] core0/mem_data_out[35]
+ core0/mem_data_out[36] core0/mem_data_out[37] core0/mem_data_out[38] core0/mem_data_out[39]
+ core0/mem_data_out[3] core0/mem_data_out[40] core0/mem_data_out[41] core0/mem_data_out[42]
+ core0/mem_data_out[43] core0/mem_data_out[44] core0/mem_data_out[45] core0/mem_data_out[46]
+ core0/mem_data_out[47] core0/mem_data_out[48] core0/mem_data_out[49] core0/mem_data_out[4]
+ core0/mem_data_out[50] core0/mem_data_out[51] core0/mem_data_out[52] core0/mem_data_out[53]
+ core0/mem_data_out[54] core0/mem_data_out[55] core0/mem_data_out[56] core0/mem_data_out[57]
+ core0/mem_data_out[58] core0/mem_data_out[59] core0/mem_data_out[5] core0/mem_data_out[60]
+ core0/mem_data_out[61] core0/mem_data_out[62] core0/mem_data_out[63] core0/mem_data_out[64]
+ core0/mem_data_out[65] core0/mem_data_out[66] core0/mem_data_out[67] core0/mem_data_out[68]
+ core0/mem_data_out[69] core0/mem_data_out[6] core0/mem_data_out[70] core0/mem_data_out[71]
+ core0/mem_data_out[72] core0/mem_data_out[73] core0/mem_data_out[74] core0/mem_data_out[75]
+ core0/mem_data_out[76] core0/mem_data_out[77] core0/mem_data_out[78] core0/mem_data_out[79]
+ core0/mem_data_out[7] core0/mem_data_out[80] core0/mem_data_out[81] core0/mem_data_out[82]
+ core0/mem_data_out[83] core0/mem_data_out[84] core0/mem_data_out[85] core0/mem_data_out[86]
+ core0/mem_data_out[87] core0/mem_data_out[88] core0/mem_data_out[89] core0/mem_data_out[8]
+ core0/mem_data_out[90] core0/mem_data_out[91] core0/mem_data_out[92] core0/mem_data_out[93]
+ core0/mem_data_out[94] core0/mem_data_out[95] core0/mem_data_out[96] core0/mem_data_out[97]
+ core0/mem_data_out[98] core0/mem_data_out[99] core0/mem_data_out[9] core0/read_interactive_ready
+ core0/read_interactive_req core0/read_interactive_value[0] core0/read_interactive_value[10]
+ core0/read_interactive_value[11] core0/read_interactive_value[12] core0/read_interactive_value[13]
+ core0/read_interactive_value[14] core0/read_interactive_value[15] core0/read_interactive_value[16]
+ core0/read_interactive_value[17] core0/read_interactive_value[18] core0/read_interactive_value[19]
+ core0/read_interactive_value[1] core0/read_interactive_value[20] core0/read_interactive_value[21]
+ core0/read_interactive_value[22] core0/read_interactive_value[23] core0/read_interactive_value[24]
+ core0/read_interactive_value[25] core0/read_interactive_value[26] core0/read_interactive_value[27]
+ core0/read_interactive_value[28] core0/read_interactive_value[29] core0/read_interactive_value[2]
+ core0/read_interactive_value[30] core0/read_interactive_value[31] core0/read_interactive_value[3]
+ core0/read_interactive_value[4] core0/read_interactive_value[5] core0/read_interactive_value[6]
+ core0/read_interactive_value[7] core0/read_interactive_value[8] core0/read_interactive_value[9]
+ core0/rst vccd1 vssd1 core
Xcustom_sram custom_sram/a[0] custom_sram/a[10] custom_sram/a[11] custom_sram/a[12]
+ custom_sram/a[13] custom_sram/a[14] custom_sram/a[15] custom_sram/a[16] custom_sram/a[17]
+ custom_sram/a[18] custom_sram/a[19] custom_sram/a[1] custom_sram/a[2] custom_sram/a[3]
+ custom_sram/a[4] custom_sram/a[5] custom_sram/a[6] custom_sram/a[7] custom_sram/a[8]
+ custom_sram/a[9] core0/clk custom_sram/csb0_to_sram custom_sram/d[0] custom_sram/d[10]
+ custom_sram/d[11] custom_sram/d[12] custom_sram/d[13] custom_sram/d[14] custom_sram/d[15]
+ custom_sram/d[16] custom_sram/d[17] custom_sram/d[18] custom_sram/d[19] custom_sram/d[1]
+ custom_sram/d[20] custom_sram/d[21] custom_sram/d[22] custom_sram/d[23] custom_sram/d[24]
+ custom_sram/d[25] custom_sram/d[26] custom_sram/d[27] custom_sram/d[28] custom_sram/d[29]
+ custom_sram/d[2] custom_sram/d[30] custom_sram/d[31] custom_sram/d[3] custom_sram/d[4]
+ custom_sram/d[5] custom_sram/d[6] custom_sram/d[7] custom_sram/d[8] custom_sram/d[9]
+ custom_sram/q[0] custom_sram/q[10] custom_sram/q[11] custom_sram/q[12] custom_sram/q[13]
+ custom_sram/q[14] custom_sram/q[15] custom_sram/q[16] custom_sram/q[17] custom_sram/q[18]
+ custom_sram/q[19] custom_sram/q[1] custom_sram/q[20] custom_sram/q[21] custom_sram/q[22]
+ custom_sram/q[23] custom_sram/q[24] custom_sram/q[25] custom_sram/q[26] custom_sram/q[27]
+ custom_sram/q[28] custom_sram/q[29] custom_sram/q[2] custom_sram/q[30] custom_sram/q[31]
+ custom_sram/q[3] custom_sram/q[4] custom_sram/q[5] custom_sram/q[6] custom_sram/q[7]
+ custom_sram/q[8] custom_sram/q[9] custom_sram/spare_wen0_to_sram vccd1 vssd1 custom_sram/we
+ custom_sram
.ends

