VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO io_input_arbiter
  CLASS BLOCK ;
  FOREIGN io_input_arbiter ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 75.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END clk
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 13.640 75.000 14.240 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 71.000 47.290 75.000 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 31.320 75.000 31.920 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 71.000 62.470 75.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 36.760 75.000 37.360 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 48.320 75.000 48.920 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 71.000 22.450 75.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 71.000 27.510 75.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 71.000 32.570 75.000 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END data_out[9]
  PIN is_ready_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 71.000 2.670 75.000 ;
    END
  END is_ready_core0
  PIN read_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 71.000 7.270 75.000 ;
    END
  END read_enable
  PIN read_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 71.000 17.390 75.000 ;
    END
  END read_value[0]
  PIN read_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END read_value[10]
  PIN read_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 19.760 75.000 20.360 ;
    END
  END read_value[11]
  PIN read_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END read_value[12]
  PIN read_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 25.200 75.000 25.800 ;
    END
  END read_value[13]
  PIN read_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 71.000 52.350 75.000 ;
    END
  END read_value[14]
  PIN read_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END read_value[15]
  PIN read_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END read_value[16]
  PIN read_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 71.000 57.410 75.000 ;
    END
  END read_value[17]
  PIN read_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END read_value[18]
  PIN read_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 71.000 67.530 75.000 ;
    END
  END read_value[19]
  PIN read_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END read_value[1]
  PIN read_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END read_value[20]
  PIN read_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END read_value[21]
  PIN read_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END read_value[22]
  PIN read_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 42.880 75.000 43.480 ;
    END
  END read_value[23]
  PIN read_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END read_value[24]
  PIN read_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 54.440 75.000 55.040 ;
    END
  END read_value[25]
  PIN read_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 59.880 75.000 60.480 ;
    END
  END read_value[26]
  PIN read_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 66.000 75.000 66.600 ;
    END
  END read_value[27]
  PIN read_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END read_value[28]
  PIN read_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END read_value[29]
  PIN read_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END read_value[2]
  PIN read_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 71.000 72.590 75.000 ;
    END
  END read_value[30]
  PIN read_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 71.440 75.000 72.040 ;
    END
  END read_value[31]
  PIN read_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 2.760 75.000 3.360 ;
    END
  END read_value[3]
  PIN read_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 8.200 75.000 8.800 ;
    END
  END read_value[4]
  PIN read_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END read_value[5]
  PIN read_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 71.000 37.630 75.000 ;
    END
  END read_value[6]
  PIN read_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END read_value[7]
  PIN read_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END read_value[8]
  PIN read_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 71.000 42.230 75.000 ;
    END
  END read_value[9]
  PIN req_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 71.000 12.330 75.000 ;
    END
  END req_core0
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.380 10.640 16.980 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.700 10.640 38.300 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.020 10.640 59.620 62.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.040 10.640 27.640 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.360 10.640 48.960 62.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 3.145 70.235 62.645 ;
      LAYER met1 ;
        RECT 1.450 3.100 73.070 62.800 ;
      LAYER met2 ;
        RECT 1.480 70.720 2.110 72.605 ;
        RECT 2.950 70.720 6.710 72.605 ;
        RECT 7.550 70.720 11.770 72.605 ;
        RECT 12.610 70.720 16.830 72.605 ;
        RECT 17.670 70.720 21.890 72.605 ;
        RECT 22.730 70.720 26.950 72.605 ;
        RECT 27.790 70.720 32.010 72.605 ;
        RECT 32.850 70.720 37.070 72.605 ;
        RECT 37.910 70.720 41.670 72.605 ;
        RECT 42.510 70.720 46.730 72.605 ;
        RECT 47.570 70.720 51.790 72.605 ;
        RECT 52.630 70.720 56.850 72.605 ;
        RECT 57.690 70.720 61.910 72.605 ;
        RECT 62.750 70.720 66.970 72.605 ;
        RECT 67.810 70.720 72.030 72.605 ;
        RECT 72.870 70.720 73.040 72.605 ;
        RECT 1.480 4.280 73.040 70.720 ;
        RECT 2.030 1.515 4.410 4.280 ;
        RECT 5.250 1.515 7.630 4.280 ;
        RECT 8.470 1.515 11.310 4.280 ;
        RECT 12.150 1.515 14.530 4.280 ;
        RECT 15.370 1.515 18.210 4.280 ;
        RECT 19.050 1.515 21.430 4.280 ;
        RECT 22.270 1.515 24.650 4.280 ;
        RECT 25.490 1.515 28.330 4.280 ;
        RECT 29.170 1.515 31.550 4.280 ;
        RECT 32.390 1.515 35.230 4.280 ;
        RECT 36.070 1.515 38.450 4.280 ;
        RECT 39.290 1.515 41.670 4.280 ;
        RECT 42.510 1.515 45.350 4.280 ;
        RECT 46.190 1.515 48.570 4.280 ;
        RECT 49.410 1.515 52.250 4.280 ;
        RECT 53.090 1.515 55.470 4.280 ;
        RECT 56.310 1.515 58.690 4.280 ;
        RECT 59.530 1.515 62.370 4.280 ;
        RECT 63.210 1.515 65.590 4.280 ;
        RECT 66.430 1.515 69.270 4.280 ;
        RECT 70.110 1.515 72.490 4.280 ;
      LAYER met3 ;
        RECT 4.400 72.440 71.000 72.585 ;
        RECT 4.400 71.720 70.600 72.440 ;
        RECT 4.000 71.040 70.600 71.720 ;
        RECT 4.000 69.040 71.000 71.040 ;
        RECT 4.400 67.640 71.000 69.040 ;
        RECT 4.000 67.000 71.000 67.640 ;
        RECT 4.000 65.600 70.600 67.000 ;
        RECT 4.000 64.960 71.000 65.600 ;
        RECT 4.400 63.560 71.000 64.960 ;
        RECT 4.000 60.880 71.000 63.560 ;
        RECT 4.400 59.480 70.600 60.880 ;
        RECT 4.000 57.480 71.000 59.480 ;
        RECT 4.400 56.080 71.000 57.480 ;
        RECT 4.000 55.440 71.000 56.080 ;
        RECT 4.000 54.040 70.600 55.440 ;
        RECT 4.000 53.400 71.000 54.040 ;
        RECT 4.400 52.000 71.000 53.400 ;
        RECT 4.000 49.320 71.000 52.000 ;
        RECT 4.400 47.920 70.600 49.320 ;
        RECT 4.000 45.240 71.000 47.920 ;
        RECT 4.400 43.880 71.000 45.240 ;
        RECT 4.400 43.840 70.600 43.880 ;
        RECT 4.000 42.480 70.600 43.840 ;
        RECT 4.000 41.160 71.000 42.480 ;
        RECT 4.400 39.760 71.000 41.160 ;
        RECT 4.000 37.760 71.000 39.760 ;
        RECT 4.400 36.360 70.600 37.760 ;
        RECT 4.000 33.680 71.000 36.360 ;
        RECT 4.400 32.320 71.000 33.680 ;
        RECT 4.400 32.280 70.600 32.320 ;
        RECT 4.000 30.920 70.600 32.280 ;
        RECT 4.000 29.600 71.000 30.920 ;
        RECT 4.400 28.200 71.000 29.600 ;
        RECT 4.000 26.200 71.000 28.200 ;
        RECT 4.000 25.520 70.600 26.200 ;
        RECT 4.400 24.800 70.600 25.520 ;
        RECT 4.400 24.120 71.000 24.800 ;
        RECT 4.000 21.440 71.000 24.120 ;
        RECT 4.400 20.760 71.000 21.440 ;
        RECT 4.400 20.040 70.600 20.760 ;
        RECT 4.000 19.360 70.600 20.040 ;
        RECT 4.000 18.040 71.000 19.360 ;
        RECT 4.400 16.640 71.000 18.040 ;
        RECT 4.000 14.640 71.000 16.640 ;
        RECT 4.000 13.960 70.600 14.640 ;
        RECT 4.400 13.240 70.600 13.960 ;
        RECT 4.400 12.560 71.000 13.240 ;
        RECT 4.000 9.880 71.000 12.560 ;
        RECT 4.400 9.200 71.000 9.880 ;
        RECT 4.400 8.480 70.600 9.200 ;
        RECT 4.000 7.800 70.600 8.480 ;
        RECT 4.000 5.800 71.000 7.800 ;
        RECT 4.400 4.400 71.000 5.800 ;
        RECT 4.000 3.760 71.000 4.400 ;
        RECT 4.000 2.400 70.600 3.760 ;
        RECT 4.400 2.360 70.600 2.400 ;
        RECT 4.400 1.535 71.000 2.360 ;
  END
END io_input_arbiter
END LIBRARY

