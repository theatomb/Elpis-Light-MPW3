VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1496.000 100.190 1500.000 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 1496.000 1252.950 1500.000 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.070 1496.000 1271.350 1500.000 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 1496.000 1289.290 1500.000 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1262.800 1500.000 1263.400 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1310.400 4.000 1311.000 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.720 4.000 1327.320 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 1496.000 1307.690 1500.000 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1311.760 1500.000 1312.360 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1359.360 4.000 1359.960 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 235.320 1500.000 235.920 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1376.360 4.000 1376.960 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 1496.000 1344.490 1500.000 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1360.720 1500.000 1361.320 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1377.040 1500.000 1377.640 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.550 1496.000 1380.830 1500.000 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.680 4.000 1393.280 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.570 0.000 1420.850 4.000 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1393.360 1500.000 1393.960 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1426.000 1500.000 1426.600 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 1496.000 374.810 1500.000 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 1496.000 1435.570 1500.000 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.090 1496.000 1472.370 1500.000 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1442.320 1500.000 1442.920 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1442.320 4.000 1442.920 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1491.280 1500.000 1491.880 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1474.960 4.000 1475.560 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 1496.000 411.150 1500.000 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 1496.000 429.550 1500.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 382.200 1500.000 382.800 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 398.520 1500.000 399.120 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 431.160 1500.000 431.760 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 1496.000 191.730 1500.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 1496.000 557.890 1500.000 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 551.520 4.000 552.120 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 1496.000 612.630 1500.000 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 561.720 1500.000 562.320 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 39.480 1500.000 40.080 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 1496.000 631.030 1500.000 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 1496.000 648.970 1500.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 627.000 1500.000 627.600 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 1496.000 667.370 1500.000 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 1496.000 685.770 1500.000 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 766.400 4.000 767.000 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 659.640 1500.000 660.240 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 88.440 1500.000 89.040 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 0.000 803.070 4.000 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 1496.000 722.110 1500.000 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 708.600 1500.000 709.200 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 724.920 1500.000 725.520 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 1496.000 740.510 1500.000 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 881.320 4.000 881.920 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 898.320 4.000 898.920 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 104.760 1500.000 105.360 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 1496.000 777.310 1500.000 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 805.840 1500.000 806.440 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 838.480 1500.000 839.080 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 1496.000 795.710 1500.000 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 1496.000 813.650 1500.000 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.280 4.000 947.880 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 0.000 873.450 4.000 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 0.000 891.390 4.000 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 4.000 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 903.760 1500.000 904.360 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 0.000 979.710 4.000 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 936.400 1500.000 937.000 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 969.040 1500.000 969.640 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 0.000 997.190 4.000 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 985.360 1500.000 985.960 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 1496.000 905.190 1500.000 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1046.560 4.000 1047.160 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.710 1496.000 941.990 1500.000 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.050 1496.000 978.330 1500.000 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1018.000 1500.000 1018.600 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.880 4.000 1063.480 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.850 1496.000 1015.130 1500.000 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1079.200 4.000 1079.800 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1066.960 1500.000 1067.560 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1099.600 1500.000 1100.200 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 1496.000 301.670 1500.000 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 1496.000 1051.470 1500.000 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 1496.000 1069.870 1500.000 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.390 1496.000 1106.670 1500.000 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1148.560 1500.000 1149.160 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1164.880 1500.000 1165.480 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.730 1496.000 1143.010 1500.000 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 0.000 1102.990 4.000 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1197.520 1500.000 1198.120 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1161.480 4.000 1162.080 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 170.040 1500.000 170.640 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.550 0.000 1173.830 4.000 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.030 0.000 1191.310 4.000 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 0.000 1208.790 4.000 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.470 1496.000 1197.750 1500.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1211.120 4.000 1211.720 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.930 0.000 1244.210 4.000 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.410 0.000 1261.690 4.000 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1230.160 1500.000 1230.760 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1246.480 1500.000 1247.080 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.270 1496.000 1234.550 1500.000 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 186.360 1500.000 186.960 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 1496.000 118.590 1500.000 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 316.920 1500.000 317.520 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 414.840 1500.000 415.440 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 1496.000 594.230 1500.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 496.440 1500.000 497.040 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 545.400 1500.000 546.000 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 578.040 1500.000 578.640 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 55.800 1500.000 56.400 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 1496.000 228.530 1500.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 137.400 1500.000 138.000 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 202.680 1500.000 203.280 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 1496.000 45.450 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 7.520 1500.000 8.120 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 1496.000 82.250 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 1496.000 63.850 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 1496.000 136.990 1500.000 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 251.640 1500.000 252.240 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 284.280 1500.000 284.880 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 349.560 1500.000 350.160 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 1496.000 466.350 1500.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 23.160 1500.000 23.760 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 1496.000 320.070 1500.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 219.000 1500.000 219.600 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 1496.000 155.390 1500.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1244.440 4.000 1245.040 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 0.000 1314.590 4.000 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1260.760 4.000 1261.360 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1277.080 4.000 1277.680 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1279.120 1500.000 1279.720 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1295.440 1500.000 1296.040 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.040 4.000 1343.640 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.250 0.000 1332.530 4.000 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1328.080 1500.000 1328.680 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.810 1496.000 1326.090 1500.000 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 1496.000 356.410 1500.000 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1344.400 1500.000 1345.000 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 0.000 1350.010 4.000 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.150 1496.000 1362.430 1500.000 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.670 0.000 1367.950 4.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.950 1496.000 1399.230 1500.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.000 4.000 1409.600 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.630 0.000 1402.910 4.000 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.050 0.000 1438.330 4.000 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1409.680 1500.000 1410.280 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 1496.000 1417.630 1500.000 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 1496.000 393.210 1500.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 1496.000 1453.970 1500.000 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.470 0.000 1473.750 4.000 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1425.320 4.000 1425.920 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1458.640 1500.000 1459.240 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1474.960 1500.000 1475.560 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 1496.000 1490.770 1500.000 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.280 4.000 1491.880 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 333.240 1500.000 333.840 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 365.880 1500.000 366.480 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 1496.000 447.950 1500.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 1496.000 484.290 1500.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 1496.000 521.090 1500.000 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 1496.000 539.490 1500.000 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 463.800 1500.000 464.400 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 512.760 1500.000 513.360 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 72.120 1500.000 72.720 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.120 4.000 667.720 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 1496.000 704.170 1500.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 643.320 1500.000 643.920 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 675.960 1500.000 676.560 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 692.280 1500.000 692.880 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 0.000 820.550 4.000 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 741.240 1500.000 741.840 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.680 4.000 849.280 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.630 1496.000 758.910 1500.000 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 757.560 1500.000 758.160 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 773.200 1500.000 773.800 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 789.520 1500.000 790.120 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 1496.000 246.470 1500.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 822.160 1500.000 822.760 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 854.800 1500.000 855.400 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 871.120 1500.000 871.720 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 1496.000 832.050 1500.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.280 4.000 964.880 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 0.000 908.870 4.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 0.000 926.350 4.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 1496.000 850.450 1500.000 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 887.440 1500.000 888.040 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 0.000 961.770 4.000 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 920.080 1500.000 920.680 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.570 1496.000 868.850 1500.000 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 952.720 1500.000 953.320 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 1496.000 886.790 1500.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 0.000 1032.610 4.000 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1001.680 1500.000 1002.280 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 1496.000 264.870 1500.000 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.310 1496.000 923.590 1500.000 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 0.000 1067.570 4.000 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 1496.000 959.930 1500.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 1496.000 996.730 1500.000 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1034.320 1500.000 1034.920 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1050.640 1500.000 1051.240 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 1496.000 1033.530 1500.000 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1083.280 1500.000 1083.880 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1095.520 4.000 1096.120 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1115.920 1500.000 1116.520 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.990 1496.000 1088.270 1500.000 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1132.240 1500.000 1132.840 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 1496.000 1124.610 1500.000 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1112.520 4.000 1113.120 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1181.200 1500.000 1181.800 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.840 4.000 1129.440 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.160 4.000 1145.760 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.610 0.000 1155.890 4.000 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1178.480 4.000 1179.080 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.130 1496.000 1161.410 1500.000 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.530 1496.000 1179.810 1500.000 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.800 4.000 1195.400 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.450 0.000 1226.730 4.000 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1213.840 1500.000 1214.440 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.350 0.000 1279.630 4.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.870 1496.000 1216.150 1500.000 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.830 0.000 1297.110 4.000 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 1496.000 9.110 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 1496.000 27.050 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 1496.000 173.330 1500.000 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 267.960 1500.000 268.560 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 300.600 1500.000 301.200 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 1496.000 502.690 1500.000 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 447.480 1500.000 448.080 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 1496.000 575.830 1500.000 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 480.120 1500.000 480.720 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 529.080 1500.000 529.680 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 634.480 4.000 635.080 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 594.360 1500.000 594.960 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 1496.000 210.130 1500.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 610.680 1500.000 611.280 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 121.080 1500.000 121.680 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 1496.000 283.270 1500.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 153.720 1500.000 154.320 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 1496.000 338.010 1500.000 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1494.855 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.915 1488.080 ;
      LAYER met2 ;
        RECT 6.600 1495.720 8.550 1496.410 ;
        RECT 9.390 1495.720 26.490 1496.410 ;
        RECT 27.330 1495.720 44.890 1496.410 ;
        RECT 45.730 1495.720 63.290 1496.410 ;
        RECT 64.130 1495.720 81.690 1496.410 ;
        RECT 82.530 1495.720 99.630 1496.410 ;
        RECT 100.470 1495.720 118.030 1496.410 ;
        RECT 118.870 1495.720 136.430 1496.410 ;
        RECT 137.270 1495.720 154.830 1496.410 ;
        RECT 155.670 1495.720 172.770 1496.410 ;
        RECT 173.610 1495.720 191.170 1496.410 ;
        RECT 192.010 1495.720 209.570 1496.410 ;
        RECT 210.410 1495.720 227.970 1496.410 ;
        RECT 228.810 1495.720 245.910 1496.410 ;
        RECT 246.750 1495.720 264.310 1496.410 ;
        RECT 265.150 1495.720 282.710 1496.410 ;
        RECT 283.550 1495.720 301.110 1496.410 ;
        RECT 301.950 1495.720 319.510 1496.410 ;
        RECT 320.350 1495.720 337.450 1496.410 ;
        RECT 338.290 1495.720 355.850 1496.410 ;
        RECT 356.690 1495.720 374.250 1496.410 ;
        RECT 375.090 1495.720 392.650 1496.410 ;
        RECT 393.490 1495.720 410.590 1496.410 ;
        RECT 411.430 1495.720 428.990 1496.410 ;
        RECT 429.830 1495.720 447.390 1496.410 ;
        RECT 448.230 1495.720 465.790 1496.410 ;
        RECT 466.630 1495.720 483.730 1496.410 ;
        RECT 484.570 1495.720 502.130 1496.410 ;
        RECT 502.970 1495.720 520.530 1496.410 ;
        RECT 521.370 1495.720 538.930 1496.410 ;
        RECT 539.770 1495.720 557.330 1496.410 ;
        RECT 558.170 1495.720 575.270 1496.410 ;
        RECT 576.110 1495.720 593.670 1496.410 ;
        RECT 594.510 1495.720 612.070 1496.410 ;
        RECT 612.910 1495.720 630.470 1496.410 ;
        RECT 631.310 1495.720 648.410 1496.410 ;
        RECT 649.250 1495.720 666.810 1496.410 ;
        RECT 667.650 1495.720 685.210 1496.410 ;
        RECT 686.050 1495.720 703.610 1496.410 ;
        RECT 704.450 1495.720 721.550 1496.410 ;
        RECT 722.390 1495.720 739.950 1496.410 ;
        RECT 740.790 1495.720 758.350 1496.410 ;
        RECT 759.190 1495.720 776.750 1496.410 ;
        RECT 777.590 1495.720 795.150 1496.410 ;
        RECT 795.990 1495.720 813.090 1496.410 ;
        RECT 813.930 1495.720 831.490 1496.410 ;
        RECT 832.330 1495.720 849.890 1496.410 ;
        RECT 850.730 1495.720 868.290 1496.410 ;
        RECT 869.130 1495.720 886.230 1496.410 ;
        RECT 887.070 1495.720 904.630 1496.410 ;
        RECT 905.470 1495.720 923.030 1496.410 ;
        RECT 923.870 1495.720 941.430 1496.410 ;
        RECT 942.270 1495.720 959.370 1496.410 ;
        RECT 960.210 1495.720 977.770 1496.410 ;
        RECT 978.610 1495.720 996.170 1496.410 ;
        RECT 997.010 1495.720 1014.570 1496.410 ;
        RECT 1015.410 1495.720 1032.970 1496.410 ;
        RECT 1033.810 1495.720 1050.910 1496.410 ;
        RECT 1051.750 1495.720 1069.310 1496.410 ;
        RECT 1070.150 1495.720 1087.710 1496.410 ;
        RECT 1088.550 1495.720 1106.110 1496.410 ;
        RECT 1106.950 1495.720 1124.050 1496.410 ;
        RECT 1124.890 1495.720 1142.450 1496.410 ;
        RECT 1143.290 1495.720 1160.850 1496.410 ;
        RECT 1161.690 1495.720 1179.250 1496.410 ;
        RECT 1180.090 1495.720 1197.190 1496.410 ;
        RECT 1198.030 1495.720 1215.590 1496.410 ;
        RECT 1216.430 1495.720 1233.990 1496.410 ;
        RECT 1234.830 1495.720 1252.390 1496.410 ;
        RECT 1253.230 1495.720 1270.790 1496.410 ;
        RECT 1271.630 1495.720 1288.730 1496.410 ;
        RECT 1289.570 1495.720 1307.130 1496.410 ;
        RECT 1307.970 1495.720 1325.530 1496.410 ;
        RECT 1326.370 1495.720 1343.930 1496.410 ;
        RECT 1344.770 1495.720 1361.870 1496.410 ;
        RECT 1362.710 1495.720 1380.270 1496.410 ;
        RECT 1381.110 1495.720 1398.670 1496.410 ;
        RECT 1399.510 1495.720 1417.070 1496.410 ;
        RECT 1417.910 1495.720 1435.010 1496.410 ;
        RECT 1435.850 1495.720 1453.410 1496.410 ;
        RECT 1454.250 1495.720 1471.810 1496.410 ;
        RECT 1472.650 1495.720 1490.210 1496.410 ;
        RECT 1491.050 1495.720 1491.220 1496.410 ;
        RECT 6.600 4.280 1491.220 1495.720 ;
        RECT 6.600 3.670 8.550 4.280 ;
        RECT 9.390 3.670 26.030 4.280 ;
        RECT 26.870 3.670 43.510 4.280 ;
        RECT 44.350 3.670 61.450 4.280 ;
        RECT 62.290 3.670 78.930 4.280 ;
        RECT 79.770 3.670 96.410 4.280 ;
        RECT 97.250 3.670 114.350 4.280 ;
        RECT 115.190 3.670 131.830 4.280 ;
        RECT 132.670 3.670 149.310 4.280 ;
        RECT 150.150 3.670 167.250 4.280 ;
        RECT 168.090 3.670 184.730 4.280 ;
        RECT 185.570 3.670 202.670 4.280 ;
        RECT 203.510 3.670 220.150 4.280 ;
        RECT 220.990 3.670 237.630 4.280 ;
        RECT 238.470 3.670 255.570 4.280 ;
        RECT 256.410 3.670 273.050 4.280 ;
        RECT 273.890 3.670 290.530 4.280 ;
        RECT 291.370 3.670 308.470 4.280 ;
        RECT 309.310 3.670 325.950 4.280 ;
        RECT 326.790 3.670 343.430 4.280 ;
        RECT 344.270 3.670 361.370 4.280 ;
        RECT 362.210 3.670 378.850 4.280 ;
        RECT 379.690 3.670 396.790 4.280 ;
        RECT 397.630 3.670 414.270 4.280 ;
        RECT 415.110 3.670 431.750 4.280 ;
        RECT 432.590 3.670 449.690 4.280 ;
        RECT 450.530 3.670 467.170 4.280 ;
        RECT 468.010 3.670 484.650 4.280 ;
        RECT 485.490 3.670 502.590 4.280 ;
        RECT 503.430 3.670 520.070 4.280 ;
        RECT 520.910 3.670 537.550 4.280 ;
        RECT 538.390 3.670 555.490 4.280 ;
        RECT 556.330 3.670 572.970 4.280 ;
        RECT 573.810 3.670 590.910 4.280 ;
        RECT 591.750 3.670 608.390 4.280 ;
        RECT 609.230 3.670 625.870 4.280 ;
        RECT 626.710 3.670 643.810 4.280 ;
        RECT 644.650 3.670 661.290 4.280 ;
        RECT 662.130 3.670 678.770 4.280 ;
        RECT 679.610 3.670 696.710 4.280 ;
        RECT 697.550 3.670 714.190 4.280 ;
        RECT 715.030 3.670 731.670 4.280 ;
        RECT 732.510 3.670 749.610 4.280 ;
        RECT 750.450 3.670 767.090 4.280 ;
        RECT 767.930 3.670 785.030 4.280 ;
        RECT 785.870 3.670 802.510 4.280 ;
        RECT 803.350 3.670 819.990 4.280 ;
        RECT 820.830 3.670 837.930 4.280 ;
        RECT 838.770 3.670 855.410 4.280 ;
        RECT 856.250 3.670 872.890 4.280 ;
        RECT 873.730 3.670 890.830 4.280 ;
        RECT 891.670 3.670 908.310 4.280 ;
        RECT 909.150 3.670 925.790 4.280 ;
        RECT 926.630 3.670 943.730 4.280 ;
        RECT 944.570 3.670 961.210 4.280 ;
        RECT 962.050 3.670 979.150 4.280 ;
        RECT 979.990 3.670 996.630 4.280 ;
        RECT 997.470 3.670 1014.110 4.280 ;
        RECT 1014.950 3.670 1032.050 4.280 ;
        RECT 1032.890 3.670 1049.530 4.280 ;
        RECT 1050.370 3.670 1067.010 4.280 ;
        RECT 1067.850 3.670 1084.950 4.280 ;
        RECT 1085.790 3.670 1102.430 4.280 ;
        RECT 1103.270 3.670 1119.910 4.280 ;
        RECT 1120.750 3.670 1137.850 4.280 ;
        RECT 1138.690 3.670 1155.330 4.280 ;
        RECT 1156.170 3.670 1173.270 4.280 ;
        RECT 1174.110 3.670 1190.750 4.280 ;
        RECT 1191.590 3.670 1208.230 4.280 ;
        RECT 1209.070 3.670 1226.170 4.280 ;
        RECT 1227.010 3.670 1243.650 4.280 ;
        RECT 1244.490 3.670 1261.130 4.280 ;
        RECT 1261.970 3.670 1279.070 4.280 ;
        RECT 1279.910 3.670 1296.550 4.280 ;
        RECT 1297.390 3.670 1314.030 4.280 ;
        RECT 1314.870 3.670 1331.970 4.280 ;
        RECT 1332.810 3.670 1349.450 4.280 ;
        RECT 1350.290 3.670 1367.390 4.280 ;
        RECT 1368.230 3.670 1384.870 4.280 ;
        RECT 1385.710 3.670 1402.350 4.280 ;
        RECT 1403.190 3.670 1420.290 4.280 ;
        RECT 1421.130 3.670 1437.770 4.280 ;
        RECT 1438.610 3.670 1455.250 4.280 ;
        RECT 1456.090 3.670 1473.190 4.280 ;
        RECT 1474.030 3.670 1490.670 4.280 ;
      LAYER met3 ;
        RECT 4.400 1490.880 1495.600 1491.745 ;
        RECT 4.000 1475.960 1496.000 1490.880 ;
        RECT 4.400 1474.560 1495.600 1475.960 ;
        RECT 4.000 1459.640 1496.000 1474.560 ;
        RECT 4.400 1458.240 1495.600 1459.640 ;
        RECT 4.000 1443.320 1496.000 1458.240 ;
        RECT 4.400 1441.920 1495.600 1443.320 ;
        RECT 4.000 1427.000 1496.000 1441.920 ;
        RECT 4.000 1426.320 1495.600 1427.000 ;
        RECT 4.400 1425.600 1495.600 1426.320 ;
        RECT 4.400 1424.920 1496.000 1425.600 ;
        RECT 4.000 1410.680 1496.000 1424.920 ;
        RECT 4.000 1410.000 1495.600 1410.680 ;
        RECT 4.400 1409.280 1495.600 1410.000 ;
        RECT 4.400 1408.600 1496.000 1409.280 ;
        RECT 4.000 1394.360 1496.000 1408.600 ;
        RECT 4.000 1393.680 1495.600 1394.360 ;
        RECT 4.400 1392.960 1495.600 1393.680 ;
        RECT 4.400 1392.280 1496.000 1392.960 ;
        RECT 4.000 1378.040 1496.000 1392.280 ;
        RECT 4.000 1377.360 1495.600 1378.040 ;
        RECT 4.400 1376.640 1495.600 1377.360 ;
        RECT 4.400 1375.960 1496.000 1376.640 ;
        RECT 4.000 1361.720 1496.000 1375.960 ;
        RECT 4.000 1360.360 1495.600 1361.720 ;
        RECT 4.400 1360.320 1495.600 1360.360 ;
        RECT 4.400 1358.960 1496.000 1360.320 ;
        RECT 4.000 1345.400 1496.000 1358.960 ;
        RECT 4.000 1344.040 1495.600 1345.400 ;
        RECT 4.400 1344.000 1495.600 1344.040 ;
        RECT 4.400 1342.640 1496.000 1344.000 ;
        RECT 4.000 1329.080 1496.000 1342.640 ;
        RECT 4.000 1327.720 1495.600 1329.080 ;
        RECT 4.400 1327.680 1495.600 1327.720 ;
        RECT 4.400 1326.320 1496.000 1327.680 ;
        RECT 4.000 1312.760 1496.000 1326.320 ;
        RECT 4.000 1311.400 1495.600 1312.760 ;
        RECT 4.400 1311.360 1495.600 1311.400 ;
        RECT 4.400 1310.000 1496.000 1311.360 ;
        RECT 4.000 1296.440 1496.000 1310.000 ;
        RECT 4.000 1295.040 1495.600 1296.440 ;
        RECT 4.000 1294.400 1496.000 1295.040 ;
        RECT 4.400 1293.000 1496.000 1294.400 ;
        RECT 4.000 1280.120 1496.000 1293.000 ;
        RECT 4.000 1278.720 1495.600 1280.120 ;
        RECT 4.000 1278.080 1496.000 1278.720 ;
        RECT 4.400 1276.680 1496.000 1278.080 ;
        RECT 4.000 1263.800 1496.000 1276.680 ;
        RECT 4.000 1262.400 1495.600 1263.800 ;
        RECT 4.000 1261.760 1496.000 1262.400 ;
        RECT 4.400 1260.360 1496.000 1261.760 ;
        RECT 4.000 1247.480 1496.000 1260.360 ;
        RECT 4.000 1246.080 1495.600 1247.480 ;
        RECT 4.000 1245.440 1496.000 1246.080 ;
        RECT 4.400 1244.040 1496.000 1245.440 ;
        RECT 4.000 1231.160 1496.000 1244.040 ;
        RECT 4.000 1229.760 1495.600 1231.160 ;
        RECT 4.000 1228.440 1496.000 1229.760 ;
        RECT 4.400 1227.040 1496.000 1228.440 ;
        RECT 4.000 1214.840 1496.000 1227.040 ;
        RECT 4.000 1213.440 1495.600 1214.840 ;
        RECT 4.000 1212.120 1496.000 1213.440 ;
        RECT 4.400 1210.720 1496.000 1212.120 ;
        RECT 4.000 1198.520 1496.000 1210.720 ;
        RECT 4.000 1197.120 1495.600 1198.520 ;
        RECT 4.000 1195.800 1496.000 1197.120 ;
        RECT 4.400 1194.400 1496.000 1195.800 ;
        RECT 4.000 1182.200 1496.000 1194.400 ;
        RECT 4.000 1180.800 1495.600 1182.200 ;
        RECT 4.000 1179.480 1496.000 1180.800 ;
        RECT 4.400 1178.080 1496.000 1179.480 ;
        RECT 4.000 1165.880 1496.000 1178.080 ;
        RECT 4.000 1164.480 1495.600 1165.880 ;
        RECT 4.000 1162.480 1496.000 1164.480 ;
        RECT 4.400 1161.080 1496.000 1162.480 ;
        RECT 4.000 1149.560 1496.000 1161.080 ;
        RECT 4.000 1148.160 1495.600 1149.560 ;
        RECT 4.000 1146.160 1496.000 1148.160 ;
        RECT 4.400 1144.760 1496.000 1146.160 ;
        RECT 4.000 1133.240 1496.000 1144.760 ;
        RECT 4.000 1131.840 1495.600 1133.240 ;
        RECT 4.000 1129.840 1496.000 1131.840 ;
        RECT 4.400 1128.440 1496.000 1129.840 ;
        RECT 4.000 1116.920 1496.000 1128.440 ;
        RECT 4.000 1115.520 1495.600 1116.920 ;
        RECT 4.000 1113.520 1496.000 1115.520 ;
        RECT 4.400 1112.120 1496.000 1113.520 ;
        RECT 4.000 1100.600 1496.000 1112.120 ;
        RECT 4.000 1099.200 1495.600 1100.600 ;
        RECT 4.000 1096.520 1496.000 1099.200 ;
        RECT 4.400 1095.120 1496.000 1096.520 ;
        RECT 4.000 1084.280 1496.000 1095.120 ;
        RECT 4.000 1082.880 1495.600 1084.280 ;
        RECT 4.000 1080.200 1496.000 1082.880 ;
        RECT 4.400 1078.800 1496.000 1080.200 ;
        RECT 4.000 1067.960 1496.000 1078.800 ;
        RECT 4.000 1066.560 1495.600 1067.960 ;
        RECT 4.000 1063.880 1496.000 1066.560 ;
        RECT 4.400 1062.480 1496.000 1063.880 ;
        RECT 4.000 1051.640 1496.000 1062.480 ;
        RECT 4.000 1050.240 1495.600 1051.640 ;
        RECT 4.000 1047.560 1496.000 1050.240 ;
        RECT 4.400 1046.160 1496.000 1047.560 ;
        RECT 4.000 1035.320 1496.000 1046.160 ;
        RECT 4.000 1033.920 1495.600 1035.320 ;
        RECT 4.000 1030.560 1496.000 1033.920 ;
        RECT 4.400 1029.160 1496.000 1030.560 ;
        RECT 4.000 1019.000 1496.000 1029.160 ;
        RECT 4.000 1017.600 1495.600 1019.000 ;
        RECT 4.000 1014.240 1496.000 1017.600 ;
        RECT 4.400 1012.840 1496.000 1014.240 ;
        RECT 4.000 1002.680 1496.000 1012.840 ;
        RECT 4.000 1001.280 1495.600 1002.680 ;
        RECT 4.000 997.920 1496.000 1001.280 ;
        RECT 4.400 996.520 1496.000 997.920 ;
        RECT 4.000 986.360 1496.000 996.520 ;
        RECT 4.000 984.960 1495.600 986.360 ;
        RECT 4.000 981.600 1496.000 984.960 ;
        RECT 4.400 980.200 1496.000 981.600 ;
        RECT 4.000 970.040 1496.000 980.200 ;
        RECT 4.000 968.640 1495.600 970.040 ;
        RECT 4.000 965.280 1496.000 968.640 ;
        RECT 4.400 963.880 1496.000 965.280 ;
        RECT 4.000 953.720 1496.000 963.880 ;
        RECT 4.000 952.320 1495.600 953.720 ;
        RECT 4.000 948.280 1496.000 952.320 ;
        RECT 4.400 946.880 1496.000 948.280 ;
        RECT 4.000 937.400 1496.000 946.880 ;
        RECT 4.000 936.000 1495.600 937.400 ;
        RECT 4.000 931.960 1496.000 936.000 ;
        RECT 4.400 930.560 1496.000 931.960 ;
        RECT 4.000 921.080 1496.000 930.560 ;
        RECT 4.000 919.680 1495.600 921.080 ;
        RECT 4.000 915.640 1496.000 919.680 ;
        RECT 4.400 914.240 1496.000 915.640 ;
        RECT 4.000 904.760 1496.000 914.240 ;
        RECT 4.000 903.360 1495.600 904.760 ;
        RECT 4.000 899.320 1496.000 903.360 ;
        RECT 4.400 897.920 1496.000 899.320 ;
        RECT 4.000 888.440 1496.000 897.920 ;
        RECT 4.000 887.040 1495.600 888.440 ;
        RECT 4.000 882.320 1496.000 887.040 ;
        RECT 4.400 880.920 1496.000 882.320 ;
        RECT 4.000 872.120 1496.000 880.920 ;
        RECT 4.000 870.720 1495.600 872.120 ;
        RECT 4.000 866.000 1496.000 870.720 ;
        RECT 4.400 864.600 1496.000 866.000 ;
        RECT 4.000 855.800 1496.000 864.600 ;
        RECT 4.000 854.400 1495.600 855.800 ;
        RECT 4.000 849.680 1496.000 854.400 ;
        RECT 4.400 848.280 1496.000 849.680 ;
        RECT 4.000 839.480 1496.000 848.280 ;
        RECT 4.000 838.080 1495.600 839.480 ;
        RECT 4.000 833.360 1496.000 838.080 ;
        RECT 4.400 831.960 1496.000 833.360 ;
        RECT 4.000 823.160 1496.000 831.960 ;
        RECT 4.000 821.760 1495.600 823.160 ;
        RECT 4.000 816.360 1496.000 821.760 ;
        RECT 4.400 814.960 1496.000 816.360 ;
        RECT 4.000 806.840 1496.000 814.960 ;
        RECT 4.000 805.440 1495.600 806.840 ;
        RECT 4.000 800.040 1496.000 805.440 ;
        RECT 4.400 798.640 1496.000 800.040 ;
        RECT 4.000 790.520 1496.000 798.640 ;
        RECT 4.000 789.120 1495.600 790.520 ;
        RECT 4.000 783.720 1496.000 789.120 ;
        RECT 4.400 782.320 1496.000 783.720 ;
        RECT 4.000 774.200 1496.000 782.320 ;
        RECT 4.000 772.800 1495.600 774.200 ;
        RECT 4.000 767.400 1496.000 772.800 ;
        RECT 4.400 766.000 1496.000 767.400 ;
        RECT 4.000 758.560 1496.000 766.000 ;
        RECT 4.000 757.160 1495.600 758.560 ;
        RECT 4.000 750.400 1496.000 757.160 ;
        RECT 4.400 749.000 1496.000 750.400 ;
        RECT 4.000 742.240 1496.000 749.000 ;
        RECT 4.000 740.840 1495.600 742.240 ;
        RECT 4.000 734.080 1496.000 740.840 ;
        RECT 4.400 732.680 1496.000 734.080 ;
        RECT 4.000 725.920 1496.000 732.680 ;
        RECT 4.000 724.520 1495.600 725.920 ;
        RECT 4.000 717.760 1496.000 724.520 ;
        RECT 4.400 716.360 1496.000 717.760 ;
        RECT 4.000 709.600 1496.000 716.360 ;
        RECT 4.000 708.200 1495.600 709.600 ;
        RECT 4.000 701.440 1496.000 708.200 ;
        RECT 4.400 700.040 1496.000 701.440 ;
        RECT 4.000 693.280 1496.000 700.040 ;
        RECT 4.000 691.880 1495.600 693.280 ;
        RECT 4.000 684.440 1496.000 691.880 ;
        RECT 4.400 683.040 1496.000 684.440 ;
        RECT 4.000 676.960 1496.000 683.040 ;
        RECT 4.000 675.560 1495.600 676.960 ;
        RECT 4.000 668.120 1496.000 675.560 ;
        RECT 4.400 666.720 1496.000 668.120 ;
        RECT 4.000 660.640 1496.000 666.720 ;
        RECT 4.000 659.240 1495.600 660.640 ;
        RECT 4.000 651.800 1496.000 659.240 ;
        RECT 4.400 650.400 1496.000 651.800 ;
        RECT 4.000 644.320 1496.000 650.400 ;
        RECT 4.000 642.920 1495.600 644.320 ;
        RECT 4.000 635.480 1496.000 642.920 ;
        RECT 4.400 634.080 1496.000 635.480 ;
        RECT 4.000 628.000 1496.000 634.080 ;
        RECT 4.000 626.600 1495.600 628.000 ;
        RECT 4.000 618.480 1496.000 626.600 ;
        RECT 4.400 617.080 1496.000 618.480 ;
        RECT 4.000 611.680 1496.000 617.080 ;
        RECT 4.000 610.280 1495.600 611.680 ;
        RECT 4.000 602.160 1496.000 610.280 ;
        RECT 4.400 600.760 1496.000 602.160 ;
        RECT 4.000 595.360 1496.000 600.760 ;
        RECT 4.000 593.960 1495.600 595.360 ;
        RECT 4.000 585.840 1496.000 593.960 ;
        RECT 4.400 584.440 1496.000 585.840 ;
        RECT 4.000 579.040 1496.000 584.440 ;
        RECT 4.000 577.640 1495.600 579.040 ;
        RECT 4.000 569.520 1496.000 577.640 ;
        RECT 4.400 568.120 1496.000 569.520 ;
        RECT 4.000 562.720 1496.000 568.120 ;
        RECT 4.000 561.320 1495.600 562.720 ;
        RECT 4.000 552.520 1496.000 561.320 ;
        RECT 4.400 551.120 1496.000 552.520 ;
        RECT 4.000 546.400 1496.000 551.120 ;
        RECT 4.000 545.000 1495.600 546.400 ;
        RECT 4.000 536.200 1496.000 545.000 ;
        RECT 4.400 534.800 1496.000 536.200 ;
        RECT 4.000 530.080 1496.000 534.800 ;
        RECT 4.000 528.680 1495.600 530.080 ;
        RECT 4.000 519.880 1496.000 528.680 ;
        RECT 4.400 518.480 1496.000 519.880 ;
        RECT 4.000 513.760 1496.000 518.480 ;
        RECT 4.000 512.360 1495.600 513.760 ;
        RECT 4.000 503.560 1496.000 512.360 ;
        RECT 4.400 502.160 1496.000 503.560 ;
        RECT 4.000 497.440 1496.000 502.160 ;
        RECT 4.000 496.040 1495.600 497.440 ;
        RECT 4.000 487.240 1496.000 496.040 ;
        RECT 4.400 485.840 1496.000 487.240 ;
        RECT 4.000 481.120 1496.000 485.840 ;
        RECT 4.000 479.720 1495.600 481.120 ;
        RECT 4.000 470.240 1496.000 479.720 ;
        RECT 4.400 468.840 1496.000 470.240 ;
        RECT 4.000 464.800 1496.000 468.840 ;
        RECT 4.000 463.400 1495.600 464.800 ;
        RECT 4.000 453.920 1496.000 463.400 ;
        RECT 4.400 452.520 1496.000 453.920 ;
        RECT 4.000 448.480 1496.000 452.520 ;
        RECT 4.000 447.080 1495.600 448.480 ;
        RECT 4.000 437.600 1496.000 447.080 ;
        RECT 4.400 436.200 1496.000 437.600 ;
        RECT 4.000 432.160 1496.000 436.200 ;
        RECT 4.000 430.760 1495.600 432.160 ;
        RECT 4.000 421.280 1496.000 430.760 ;
        RECT 4.400 419.880 1496.000 421.280 ;
        RECT 4.000 415.840 1496.000 419.880 ;
        RECT 4.000 414.440 1495.600 415.840 ;
        RECT 4.000 404.280 1496.000 414.440 ;
        RECT 4.400 402.880 1496.000 404.280 ;
        RECT 4.000 399.520 1496.000 402.880 ;
        RECT 4.000 398.120 1495.600 399.520 ;
        RECT 4.000 387.960 1496.000 398.120 ;
        RECT 4.400 386.560 1496.000 387.960 ;
        RECT 4.000 383.200 1496.000 386.560 ;
        RECT 4.000 381.800 1495.600 383.200 ;
        RECT 4.000 371.640 1496.000 381.800 ;
        RECT 4.400 370.240 1496.000 371.640 ;
        RECT 4.000 366.880 1496.000 370.240 ;
        RECT 4.000 365.480 1495.600 366.880 ;
        RECT 4.000 355.320 1496.000 365.480 ;
        RECT 4.400 353.920 1496.000 355.320 ;
        RECT 4.000 350.560 1496.000 353.920 ;
        RECT 4.000 349.160 1495.600 350.560 ;
        RECT 4.000 338.320 1496.000 349.160 ;
        RECT 4.400 336.920 1496.000 338.320 ;
        RECT 4.000 334.240 1496.000 336.920 ;
        RECT 4.000 332.840 1495.600 334.240 ;
        RECT 4.000 322.000 1496.000 332.840 ;
        RECT 4.400 320.600 1496.000 322.000 ;
        RECT 4.000 317.920 1496.000 320.600 ;
        RECT 4.000 316.520 1495.600 317.920 ;
        RECT 4.000 305.680 1496.000 316.520 ;
        RECT 4.400 304.280 1496.000 305.680 ;
        RECT 4.000 301.600 1496.000 304.280 ;
        RECT 4.000 300.200 1495.600 301.600 ;
        RECT 4.000 289.360 1496.000 300.200 ;
        RECT 4.400 287.960 1496.000 289.360 ;
        RECT 4.000 285.280 1496.000 287.960 ;
        RECT 4.000 283.880 1495.600 285.280 ;
        RECT 4.000 272.360 1496.000 283.880 ;
        RECT 4.400 270.960 1496.000 272.360 ;
        RECT 4.000 268.960 1496.000 270.960 ;
        RECT 4.000 267.560 1495.600 268.960 ;
        RECT 4.000 256.040 1496.000 267.560 ;
        RECT 4.400 254.640 1496.000 256.040 ;
        RECT 4.000 252.640 1496.000 254.640 ;
        RECT 4.000 251.240 1495.600 252.640 ;
        RECT 4.000 239.720 1496.000 251.240 ;
        RECT 4.400 238.320 1496.000 239.720 ;
        RECT 4.000 236.320 1496.000 238.320 ;
        RECT 4.000 234.920 1495.600 236.320 ;
        RECT 4.000 223.400 1496.000 234.920 ;
        RECT 4.400 222.000 1496.000 223.400 ;
        RECT 4.000 220.000 1496.000 222.000 ;
        RECT 4.000 218.600 1495.600 220.000 ;
        RECT 4.000 206.400 1496.000 218.600 ;
        RECT 4.400 205.000 1496.000 206.400 ;
        RECT 4.000 203.680 1496.000 205.000 ;
        RECT 4.000 202.280 1495.600 203.680 ;
        RECT 4.000 190.080 1496.000 202.280 ;
        RECT 4.400 188.680 1496.000 190.080 ;
        RECT 4.000 187.360 1496.000 188.680 ;
        RECT 4.000 185.960 1495.600 187.360 ;
        RECT 4.000 173.760 1496.000 185.960 ;
        RECT 4.400 172.360 1496.000 173.760 ;
        RECT 4.000 171.040 1496.000 172.360 ;
        RECT 4.000 169.640 1495.600 171.040 ;
        RECT 4.000 157.440 1496.000 169.640 ;
        RECT 4.400 156.040 1496.000 157.440 ;
        RECT 4.000 154.720 1496.000 156.040 ;
        RECT 4.000 153.320 1495.600 154.720 ;
        RECT 4.000 140.440 1496.000 153.320 ;
        RECT 4.400 139.040 1496.000 140.440 ;
        RECT 4.000 138.400 1496.000 139.040 ;
        RECT 4.000 137.000 1495.600 138.400 ;
        RECT 4.000 124.120 1496.000 137.000 ;
        RECT 4.400 122.720 1496.000 124.120 ;
        RECT 4.000 122.080 1496.000 122.720 ;
        RECT 4.000 120.680 1495.600 122.080 ;
        RECT 4.000 107.800 1496.000 120.680 ;
        RECT 4.400 106.400 1496.000 107.800 ;
        RECT 4.000 105.760 1496.000 106.400 ;
        RECT 4.000 104.360 1495.600 105.760 ;
        RECT 4.000 91.480 1496.000 104.360 ;
        RECT 4.400 90.080 1496.000 91.480 ;
        RECT 4.000 89.440 1496.000 90.080 ;
        RECT 4.000 88.040 1495.600 89.440 ;
        RECT 4.000 74.480 1496.000 88.040 ;
        RECT 4.400 73.120 1496.000 74.480 ;
        RECT 4.400 73.080 1495.600 73.120 ;
        RECT 4.000 71.720 1495.600 73.080 ;
        RECT 4.000 58.160 1496.000 71.720 ;
        RECT 4.400 56.800 1496.000 58.160 ;
        RECT 4.400 56.760 1495.600 56.800 ;
        RECT 4.000 55.400 1495.600 56.760 ;
        RECT 4.000 41.840 1496.000 55.400 ;
        RECT 4.400 40.480 1496.000 41.840 ;
        RECT 4.400 40.440 1495.600 40.480 ;
        RECT 4.000 39.080 1495.600 40.440 ;
        RECT 4.000 25.520 1496.000 39.080 ;
        RECT 4.400 24.160 1496.000 25.520 ;
        RECT 4.400 24.120 1495.600 24.160 ;
        RECT 4.000 22.760 1495.600 24.120 ;
        RECT 4.000 9.200 1496.000 22.760 ;
        RECT 4.400 8.520 1496.000 9.200 ;
        RECT 4.400 7.800 1495.600 8.520 ;
        RECT 4.000 7.655 1495.600 7.800 ;
      LAYER met4 ;
        RECT 100.575 11.735 174.240 1485.625 ;
        RECT 176.640 11.735 251.040 1485.625 ;
        RECT 253.440 11.735 327.840 1485.625 ;
        RECT 330.240 11.735 404.640 1485.625 ;
        RECT 407.040 11.735 481.440 1485.625 ;
        RECT 483.840 11.735 558.240 1485.625 ;
        RECT 560.640 11.735 635.040 1485.625 ;
        RECT 637.440 11.735 711.840 1485.625 ;
        RECT 714.240 11.735 788.640 1485.625 ;
        RECT 791.040 11.735 865.440 1485.625 ;
        RECT 867.840 11.735 942.240 1485.625 ;
        RECT 944.640 11.735 1019.040 1485.625 ;
        RECT 1021.440 11.735 1095.840 1485.625 ;
        RECT 1098.240 11.735 1172.640 1485.625 ;
        RECT 1175.040 11.735 1200.305 1485.625 ;
  END
END core
END LIBRARY

