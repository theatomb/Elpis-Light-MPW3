VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO custom_sram
  CLASS BLOCK ;
  FOREIGN custom_sram ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 1500.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 862.280 1800.000 862.880 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 1496.000 642.990 1500.000 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1087.360 1800.000 1087.960 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1162.160 1800.000 1162.760 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1496.000 900.130 1500.000 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 0.000 1242.830 4.000 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 1496.000 1242.830 1500.000 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 187.040 1800.000 187.640 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 1496.000 214.270 1500.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 412.120 1800.000 412.720 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 486.920 1800.000 487.520 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 637.200 1800.000 637.800 ;
    END
  END a[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END clk
  PIN csb0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END csb0_to_sram
  PIN d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END d[0]
  PIN d[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END d[10]
  PIN d[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 787.480 1800.000 788.080 ;
    END
  END d[11]
  PIN d[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 937.080 1800.000 937.680 ;
    END
  END d[12]
  PIN d[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1011.880 1800.000 1012.480 ;
    END
  END d[13]
  PIN d[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 0.000 1071.710 4.000 ;
    END
  END d[14]
  PIN d[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 0.000 1157.270 4.000 ;
    END
  END d[15]
  PIN d[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 1496.000 728.550 1500.000 ;
    END
  END d[16]
  PIN d[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 1496.000 985.690 1500.000 ;
    END
  END d[17]
  PIN d[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END d[18]
  PIN d[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1236.960 1800.000 1237.560 ;
    END
  END d[19]
  PIN d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 37.440 1800.000 38.040 ;
    END
  END d[1]
  PIN d[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1312.440 1800.000 1313.040 ;
    END
  END d[20]
  PIN d[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.160 4.000 1009.760 ;
    END
  END d[21]
  PIN d[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 0.000 1499.970 4.000 ;
    END
  END d[22]
  PIN d[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.570 1496.000 1328.850 1500.000 ;
    END
  END d[23]
  PIN d[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 1496.000 1499.970 1500.000 ;
    END
  END d[24]
  PIN d[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.710 1496.000 1585.990 1500.000 ;
    END
  END d[25]
  PIN d[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.680 4.000 1240.280 ;
    END
  END d[26]
  PIN d[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 1496.000 1671.550 1500.000 ;
    END
  END d[27]
  PIN d[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1387.240 1800.000 1387.840 ;
    END
  END d[28]
  PIN d[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 0.000 1671.550 4.000 ;
    END
  END d[29]
  PIN d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 1496.000 128.710 1500.000 ;
    END
  END d[2]
  PIN d[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1355.280 4.000 1355.880 ;
    END
  END d[30]
  PIN d[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1470.880 4.000 1471.480 ;
    END
  END d[31]
  PIN d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 261.840 1800.000 262.440 ;
    END
  END d[3]
  PIN d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 1496.000 300.290 1500.000 ;
    END
  END d[4]
  PIN d[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END d[5]
  PIN d[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END d[6]
  PIN d[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 562.400 1800.000 563.000 ;
    END
  END d[7]
  PIN d[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 1496.000 385.850 1500.000 ;
    END
  END d[8]
  PIN d[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 1496.000 471.410 1500.000 ;
    END
  END d[9]
  PIN q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 1496.000 43.150 1500.000 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 712.000 1800.000 712.600 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 0.000 900.130 4.000 ;
    END
  END q[11]
  PIN q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 1496.000 557.430 1500.000 ;
    END
  END q[12]
  PIN q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END q[13]
  PIN q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END q[14]
  PIN q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.760 4.000 836.360 ;
    END
  END q[15]
  PIN q[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 1496.000 814.570 1500.000 ;
    END
  END q[16]
  PIN q[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 1496.000 1071.710 1500.000 ;
    END
  END q[17]
  PIN q[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 1496.000 1157.270 1500.000 ;
    END
  END q[18]
  PIN q[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.570 0.000 1328.850 4.000 ;
    END
  END q[19]
  PIN q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 112.240 1800.000 112.840 ;
    END
  END q[1]
  PIN q[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 951.360 4.000 951.960 ;
    END
  END q[20]
  PIN q[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.130 0.000 1414.410 4.000 ;
    END
  END q[21]
  PIN q[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.960 4.000 1067.560 ;
    END
  END q[22]
  PIN q[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.130 1496.000 1414.410 1500.000 ;
    END
  END q[23]
  PIN q[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.760 4.000 1125.360 ;
    END
  END q[24]
  PIN q[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1181.880 4.000 1182.480 ;
    END
  END q[25]
  PIN q[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.710 0.000 1585.990 4.000 ;
    END
  END q[26]
  PIN q[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.830 1496.000 1757.110 1500.000 ;
    END
  END q[27]
  PIN q[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1297.480 4.000 1298.080 ;
    END
  END q[28]
  PIN q[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1462.040 1800.000 1462.640 ;
    END
  END q[29]
  PIN q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END q[2]
  PIN q[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1413.080 4.000 1413.680 ;
    END
  END q[30]
  PIN q[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.830 0.000 1757.110 4.000 ;
    END
  END q[31]
  PIN q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 337.320 1800.000 337.920 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END q[9]
  PIN spare_wen0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1488.080 ;
    END
  END vssd1
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END we
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1797.075 1487.925 ;
      LAYER met1 ;
        RECT 5.520 8.540 1797.135 1488.080 ;
      LAYER met2 ;
        RECT 6.990 1495.720 42.590 1496.000 ;
        RECT 43.430 1495.720 128.150 1496.000 ;
        RECT 128.990 1495.720 213.710 1496.000 ;
        RECT 214.550 1495.720 299.730 1496.000 ;
        RECT 300.570 1495.720 385.290 1496.000 ;
        RECT 386.130 1495.720 470.850 1496.000 ;
        RECT 471.690 1495.720 556.870 1496.000 ;
        RECT 557.710 1495.720 642.430 1496.000 ;
        RECT 643.270 1495.720 727.990 1496.000 ;
        RECT 728.830 1495.720 814.010 1496.000 ;
        RECT 814.850 1495.720 899.570 1496.000 ;
        RECT 900.410 1495.720 985.130 1496.000 ;
        RECT 985.970 1495.720 1071.150 1496.000 ;
        RECT 1071.990 1495.720 1156.710 1496.000 ;
        RECT 1157.550 1495.720 1242.270 1496.000 ;
        RECT 1243.110 1495.720 1328.290 1496.000 ;
        RECT 1329.130 1495.720 1413.850 1496.000 ;
        RECT 1414.690 1495.720 1499.410 1496.000 ;
        RECT 1500.250 1495.720 1585.430 1496.000 ;
        RECT 1586.270 1495.720 1670.990 1496.000 ;
        RECT 1671.830 1495.720 1756.550 1496.000 ;
        RECT 1757.390 1495.720 1792.530 1496.000 ;
        RECT 6.990 4.280 1792.530 1495.720 ;
        RECT 6.990 3.670 42.590 4.280 ;
        RECT 43.430 3.670 128.150 4.280 ;
        RECT 128.990 3.670 213.710 4.280 ;
        RECT 214.550 3.670 299.730 4.280 ;
        RECT 300.570 3.670 385.290 4.280 ;
        RECT 386.130 3.670 470.850 4.280 ;
        RECT 471.690 3.670 556.870 4.280 ;
        RECT 557.710 3.670 642.430 4.280 ;
        RECT 643.270 3.670 727.990 4.280 ;
        RECT 728.830 3.670 814.010 4.280 ;
        RECT 814.850 3.670 899.570 4.280 ;
        RECT 900.410 3.670 985.130 4.280 ;
        RECT 985.970 3.670 1071.150 4.280 ;
        RECT 1071.990 3.670 1156.710 4.280 ;
        RECT 1157.550 3.670 1242.270 4.280 ;
        RECT 1243.110 3.670 1328.290 4.280 ;
        RECT 1329.130 3.670 1413.850 4.280 ;
        RECT 1414.690 3.670 1499.410 4.280 ;
        RECT 1500.250 3.670 1585.430 4.280 ;
        RECT 1586.270 3.670 1670.990 4.280 ;
        RECT 1671.830 3.670 1756.550 4.280 ;
        RECT 1757.390 3.670 1792.530 4.280 ;
      LAYER met3 ;
        RECT 4.000 1471.880 1796.000 1488.005 ;
        RECT 4.400 1470.480 1796.000 1471.880 ;
        RECT 4.000 1463.040 1796.000 1470.480 ;
        RECT 4.000 1461.640 1795.600 1463.040 ;
        RECT 4.000 1414.080 1796.000 1461.640 ;
        RECT 4.400 1412.680 1796.000 1414.080 ;
        RECT 4.000 1388.240 1796.000 1412.680 ;
        RECT 4.000 1386.840 1795.600 1388.240 ;
        RECT 4.000 1356.280 1796.000 1386.840 ;
        RECT 4.400 1354.880 1796.000 1356.280 ;
        RECT 4.000 1313.440 1796.000 1354.880 ;
        RECT 4.000 1312.040 1795.600 1313.440 ;
        RECT 4.000 1298.480 1796.000 1312.040 ;
        RECT 4.400 1297.080 1796.000 1298.480 ;
        RECT 4.000 1240.680 1796.000 1297.080 ;
        RECT 4.400 1239.280 1796.000 1240.680 ;
        RECT 4.000 1237.960 1796.000 1239.280 ;
        RECT 4.000 1236.560 1795.600 1237.960 ;
        RECT 4.000 1182.880 1796.000 1236.560 ;
        RECT 4.400 1181.480 1796.000 1182.880 ;
        RECT 4.000 1163.160 1796.000 1181.480 ;
        RECT 4.000 1161.760 1795.600 1163.160 ;
        RECT 4.000 1125.760 1796.000 1161.760 ;
        RECT 4.400 1124.360 1796.000 1125.760 ;
        RECT 4.000 1088.360 1796.000 1124.360 ;
        RECT 4.000 1086.960 1795.600 1088.360 ;
        RECT 4.000 1067.960 1796.000 1086.960 ;
        RECT 4.400 1066.560 1796.000 1067.960 ;
        RECT 4.000 1012.880 1796.000 1066.560 ;
        RECT 4.000 1011.480 1795.600 1012.880 ;
        RECT 4.000 1010.160 1796.000 1011.480 ;
        RECT 4.400 1008.760 1796.000 1010.160 ;
        RECT 4.000 952.360 1796.000 1008.760 ;
        RECT 4.400 950.960 1796.000 952.360 ;
        RECT 4.000 938.080 1796.000 950.960 ;
        RECT 4.000 936.680 1795.600 938.080 ;
        RECT 4.000 894.560 1796.000 936.680 ;
        RECT 4.400 893.160 1796.000 894.560 ;
        RECT 4.000 863.280 1796.000 893.160 ;
        RECT 4.000 861.880 1795.600 863.280 ;
        RECT 4.000 836.760 1796.000 861.880 ;
        RECT 4.400 835.360 1796.000 836.760 ;
        RECT 4.000 788.480 1796.000 835.360 ;
        RECT 4.000 787.080 1795.600 788.480 ;
        RECT 4.000 779.640 1796.000 787.080 ;
        RECT 4.400 778.240 1796.000 779.640 ;
        RECT 4.000 721.840 1796.000 778.240 ;
        RECT 4.400 720.440 1796.000 721.840 ;
        RECT 4.000 713.000 1796.000 720.440 ;
        RECT 4.000 711.600 1795.600 713.000 ;
        RECT 4.000 664.040 1796.000 711.600 ;
        RECT 4.400 662.640 1796.000 664.040 ;
        RECT 4.000 638.200 1796.000 662.640 ;
        RECT 4.000 636.800 1795.600 638.200 ;
        RECT 4.000 606.240 1796.000 636.800 ;
        RECT 4.400 604.840 1796.000 606.240 ;
        RECT 4.000 563.400 1796.000 604.840 ;
        RECT 4.000 562.000 1795.600 563.400 ;
        RECT 4.000 548.440 1796.000 562.000 ;
        RECT 4.400 547.040 1796.000 548.440 ;
        RECT 4.000 490.640 1796.000 547.040 ;
        RECT 4.400 489.240 1796.000 490.640 ;
        RECT 4.000 487.920 1796.000 489.240 ;
        RECT 4.000 486.520 1795.600 487.920 ;
        RECT 4.000 432.840 1796.000 486.520 ;
        RECT 4.400 431.440 1796.000 432.840 ;
        RECT 4.000 413.120 1796.000 431.440 ;
        RECT 4.000 411.720 1795.600 413.120 ;
        RECT 4.000 375.720 1796.000 411.720 ;
        RECT 4.400 374.320 1796.000 375.720 ;
        RECT 4.000 338.320 1796.000 374.320 ;
        RECT 4.000 336.920 1795.600 338.320 ;
        RECT 4.000 317.920 1796.000 336.920 ;
        RECT 4.400 316.520 1796.000 317.920 ;
        RECT 4.000 262.840 1796.000 316.520 ;
        RECT 4.000 261.440 1795.600 262.840 ;
        RECT 4.000 260.120 1796.000 261.440 ;
        RECT 4.400 258.720 1796.000 260.120 ;
        RECT 4.000 202.320 1796.000 258.720 ;
        RECT 4.400 200.920 1796.000 202.320 ;
        RECT 4.000 188.040 1796.000 200.920 ;
        RECT 4.000 186.640 1795.600 188.040 ;
        RECT 4.000 144.520 1796.000 186.640 ;
        RECT 4.400 143.120 1796.000 144.520 ;
        RECT 4.000 113.240 1796.000 143.120 ;
        RECT 4.000 111.840 1795.600 113.240 ;
        RECT 4.000 86.720 1796.000 111.840 ;
        RECT 4.400 85.320 1796.000 86.720 ;
        RECT 4.000 38.440 1796.000 85.320 ;
        RECT 4.000 37.040 1795.600 38.440 ;
        RECT 4.000 29.600 1796.000 37.040 ;
        RECT 4.400 28.200 1796.000 29.600 ;
        RECT 4.000 10.715 1796.000 28.200 ;
      LAYER met4 ;
        RECT 23.295 15.135 97.440 1484.265 ;
        RECT 99.840 15.135 174.240 1484.265 ;
        RECT 176.640 15.135 251.040 1484.265 ;
        RECT 253.440 15.135 327.840 1484.265 ;
        RECT 330.240 15.135 404.640 1484.265 ;
        RECT 407.040 15.135 481.440 1484.265 ;
        RECT 483.840 15.135 558.240 1484.265 ;
        RECT 560.640 15.135 635.040 1484.265 ;
        RECT 637.440 15.135 711.840 1484.265 ;
        RECT 714.240 15.135 788.640 1484.265 ;
        RECT 791.040 15.135 865.440 1484.265 ;
        RECT 867.840 15.135 942.240 1484.265 ;
        RECT 944.640 15.135 1019.040 1484.265 ;
        RECT 1021.440 15.135 1095.840 1484.265 ;
        RECT 1098.240 15.135 1172.640 1484.265 ;
        RECT 1175.040 15.135 1249.440 1484.265 ;
        RECT 1251.840 15.135 1326.240 1484.265 ;
        RECT 1328.640 15.135 1403.040 1484.265 ;
        RECT 1405.440 15.135 1479.840 1484.265 ;
        RECT 1482.240 15.135 1556.640 1484.265 ;
        RECT 1559.040 15.135 1633.440 1484.265 ;
        RECT 1635.840 15.135 1710.240 1484.265 ;
        RECT 1712.640 15.135 1784.505 1484.265 ;
  END
END custom_sram
END LIBRARY

