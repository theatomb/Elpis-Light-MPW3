VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MEM_WB
  CLASS BLOCK ;
  FOREIGN MEM_WB ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END clk
  PIN exc_code_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 796.000 617.690 800.000 ;
    END
  END exc_code_in[0]
  PIN exc_code_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 560.360 800.000 560.960 ;
    END
  END exc_code_in[10]
  PIN exc_code_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END exc_code_in[11]
  PIN exc_code_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END exc_code_in[12]
  PIN exc_code_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END exc_code_in[13]
  PIN exc_code_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END exc_code_in[14]
  PIN exc_code_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 458.360 800.000 458.960 ;
    END
  END exc_code_in[15]
  PIN exc_code_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END exc_code_in[16]
  PIN exc_code_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END exc_code_in[17]
  PIN exc_code_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 796.000 664.610 800.000 ;
    END
  END exc_code_in[18]
  PIN exc_code_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END exc_code_in[19]
  PIN exc_code_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 287.000 800.000 287.600 ;
    END
  END exc_code_in[1]
  PIN exc_code_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 210.840 800.000 211.440 ;
    END
  END exc_code_in[20]
  PIN exc_code_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END exc_code_in[21]
  PIN exc_code_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END exc_code_in[22]
  PIN exc_code_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 216.280 800.000 216.880 ;
    END
  END exc_code_in[23]
  PIN exc_code_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END exc_code_in[24]
  PIN exc_code_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 796.000 359.170 800.000 ;
    END
  END exc_code_in[25]
  PIN exc_code_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 470.600 800.000 471.200 ;
    END
  END exc_code_in[26]
  PIN exc_code_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 330.520 800.000 331.120 ;
    END
  END exc_code_in[27]
  PIN exc_code_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 280.200 800.000 280.800 ;
    END
  END exc_code_in[28]
  PIN exc_code_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 796.000 160.450 800.000 ;
    END
  END exc_code_in[29]
  PIN exc_code_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 389.000 800.000 389.600 ;
    END
  END exc_code_in[2]
  PIN exc_code_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 796.000 647.130 800.000 ;
    END
  END exc_code_in[30]
  PIN exc_code_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END exc_code_in[31]
  PIN exc_code_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 541.320 800.000 541.920 ;
    END
  END exc_code_in[3]
  PIN exc_code_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END exc_code_in[4]
  PIN exc_code_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END exc_code_in[5]
  PIN exc_code_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END exc_code_in[6]
  PIN exc_code_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END exc_code_in[7]
  PIN exc_code_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END exc_code_in[8]
  PIN exc_code_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 796.000 595.610 800.000 ;
    END
  END exc_code_in[9]
  PIN flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 796.000 341.690 800.000 ;
    END
  END flush
  PIN io_code_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 796.000 389.530 800.000 ;
    END
  END io_code_in[0]
  PIN io_code_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END io_code_in[1]
  PIN io_code_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 796.000 634.250 800.000 ;
    END
  END io_code_in[2]
  PIN io_code_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 796.000 212.890 800.000 ;
    END
  END io_code_in[3]
  PIN io_code_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 796.000 759.370 800.000 ;
    END
  END io_code_in[4]
  PIN io_code_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END io_code_in[5]
  PIN io_code_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 796.000 354.570 800.000 ;
    END
  END io_code_in[6]
  PIN io_code_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 756.200 4.000 756.800 ;
    END
  END io_code_out[0]
  PIN io_code_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 796.000 238.650 800.000 ;
    END
  END io_code_out[1]
  PIN io_code_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 796.000 410.690 800.000 ;
    END
  END io_code_out[2]
  PIN io_code_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END io_code_out[3]
  PIN io_code_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 796.000 242.330 800.000 ;
    END
  END io_code_out[4]
  PIN io_code_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 796.000 31.650 800.000 ;
    END
  END io_code_out[5]
  PIN io_code_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 796.000 380.330 800.000 ;
    END
  END io_code_out[6]
  PIN is_ecall_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END is_ecall_in
  PIN is_flush_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 795.640 800.000 796.240 ;
    END
  END is_flush_in
  PIN is_flush_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END is_flush_out
  PIN is_hit_dtlb_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 796.000 285.570 800.000 ;
    END
  END is_hit_dtlb_in
  PIN is_hit_dtlb_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 796.000 1.290 800.000 ;
    END
  END is_hit_dtlb_out
  PIN is_hit_itlb_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END is_hit_itlb_in
  PIN is_hit_itlb_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 796.000 613.090 800.000 ;
    END
  END is_hit_itlb_out
  PIN is_iret_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END is_iret_in
  PIN is_iret_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END is_iret_out
  PIN is_mov_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END is_mov_in[0]
  PIN is_mov_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END is_mov_in[1]
  PIN is_mov_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 796.000 165.050 800.000 ;
    END
  END is_mov_out[0]
  PIN is_mov_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 796.000 203.690 800.000 ;
    END
  END is_mov_out[1]
  PIN is_read_interactive_enabled_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 465.160 800.000 465.760 ;
    END
  END is_read_interactive_enabled_in
  PIN is_read_interactive_enabled_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 796.000 221.170 800.000 ;
    END
  END is_read_interactive_enabled_out
  PIN mem_addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 796.000 182.530 800.000 ;
    END
  END mem_addr_in[0]
  PIN mem_addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END mem_addr_in[10]
  PIN mem_addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END mem_addr_in[11]
  PIN mem_addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END mem_addr_in[12]
  PIN mem_addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END mem_addr_in[13]
  PIN mem_addr_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 242.120 800.000 242.720 ;
    END
  END mem_addr_in[14]
  PIN mem_addr_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 254.360 800.000 254.960 ;
    END
  END mem_addr_in[15]
  PIN mem_addr_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END mem_addr_in[16]
  PIN mem_addr_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 477.400 800.000 478.000 ;
    END
  END mem_addr_in[17]
  PIN mem_addr_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 796.000 651.730 800.000 ;
    END
  END mem_addr_in[18]
  PIN mem_addr_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END mem_addr_in[19]
  PIN mem_addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END mem_addr_in[1]
  PIN mem_addr_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 796.000 36.250 800.000 ;
    END
  END mem_addr_in[20]
  PIN mem_addr_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END mem_addr_in[21]
  PIN mem_addr_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END mem_addr_in[22]
  PIN mem_addr_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END mem_addr_in[23]
  PIN mem_addr_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END mem_addr_in[24]
  PIN mem_addr_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END mem_addr_in[25]
  PIN mem_addr_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 261.160 800.000 261.760 ;
    END
  END mem_addr_in[26]
  PIN mem_addr_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END mem_addr_in[27]
  PIN mem_addr_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 796.000 505.450 800.000 ;
    END
  END mem_addr_in[28]
  PIN mem_addr_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END mem_addr_in[29]
  PIN mem_addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 548.120 800.000 548.720 ;
    END
  END mem_addr_in[2]
  PIN mem_addr_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 796.000 441.050 800.000 ;
    END
  END mem_addr_in[30]
  PIN mem_addr_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 796.000 716.130 800.000 ;
    END
  END mem_addr_in[31]
  PIN mem_addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END mem_addr_in[3]
  PIN mem_addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 796.000 712.450 800.000 ;
    END
  END mem_addr_in[4]
  PIN mem_addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 4.000 ;
    END
  END mem_addr_in[5]
  PIN mem_addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END mem_addr_in[6]
  PIN mem_addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 707.240 800.000 707.840 ;
    END
  END mem_addr_in[7]
  PIN mem_addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END mem_addr_in[8]
  PIN mem_addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END mem_addr_in[9]
  PIN mem_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END mem_data_in[0]
  PIN mem_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END mem_data_in[10]
  PIN mem_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END mem_data_in[11]
  PIN mem_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 796.000 324.210 800.000 ;
    END
  END mem_data_in[12]
  PIN mem_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END mem_data_in[13]
  PIN mem_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END mem_data_in[14]
  PIN mem_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 534.520 800.000 535.120 ;
    END
  END mem_data_in[15]
  PIN mem_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END mem_data_in[16]
  PIN mem_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 325.080 800.000 325.680 ;
    END
  END mem_data_in[17]
  PIN mem_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 796.000 741.890 800.000 ;
    END
  END mem_data_in[18]
  PIN mem_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END mem_data_in[19]
  PIN mem_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END mem_data_in[1]
  PIN mem_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END mem_data_in[20]
  PIN mem_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 796.000 582.730 800.000 ;
    END
  END mem_data_in[21]
  PIN mem_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 617.480 800.000 618.080 ;
    END
  END mem_data_in[22]
  PIN mem_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 700.440 800.000 701.040 ;
    END
  END mem_data_in[23]
  PIN mem_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 796.000 462.210 800.000 ;
    END
  END mem_data_in[24]
  PIN mem_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 796.000 200.010 800.000 ;
    END
  END mem_data_in[25]
  PIN mem_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 796.000 729.010 800.000 ;
    END
  END mem_data_in[26]
  PIN mem_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END mem_data_in[27]
  PIN mem_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 178.200 800.000 178.800 ;
    END
  END mem_data_in[28]
  PIN mem_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END mem_data_in[29]
  PIN mem_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 796.000 402.410 800.000 ;
    END
  END mem_data_in[2]
  PIN mem_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 796.000 510.050 800.000 ;
    END
  END mem_data_in[30]
  PIN mem_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END mem_data_in[31]
  PIN mem_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END mem_data_in[3]
  PIN mem_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END mem_data_in[4]
  PIN mem_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END mem_data_in[5]
  PIN mem_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END mem_data_in[6]
  PIN mem_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END mem_data_in[7]
  PIN mem_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END mem_data_in[8]
  PIN mem_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END mem_data_in[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 796.000 280.970 800.000 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 0.000 701.410 4.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 796.000 475.090 800.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 796.000 793.410 800.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 796.000 565.250 800.000 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 796.000 767.650 800.000 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 586.200 800.000 586.800 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 796.000 121.810 800.000 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 796.000 259.810 800.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 503.240 800.000 503.840 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 796.000 397.810 800.000 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 796.000 87.770 800.000 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 610.680 800.000 611.280 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 44.920 800.000 45.520 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 796.000 483.370 800.000 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 796.000 733.610 800.000 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 796.000 630.570 800.000 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 446.120 800.000 446.720 ;
    END
  END mem_data_out[9]
  PIN mem_to_reg_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END mem_to_reg_in
  PIN mem_to_reg_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END mem_to_reg_out
  PIN pc_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END pc_in[0]
  PIN pc_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 235.320 800.000 235.920 ;
    END
  END pc_in[10]
  PIN pc_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END pc_in[11]
  PIN pc_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 522.280 800.000 522.880 ;
    END
  END pc_in[12]
  PIN pc_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 796.000 682.090 800.000 ;
    END
  END pc_in[13]
  PIN pc_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 4.000 ;
    END
  END pc_in[14]
  PIN pc_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END pc_in[15]
  PIN pc_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END pc_in[16]
  PIN pc_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 796.000 234.050 800.000 ;
    END
  END pc_in[17]
  PIN pc_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END pc_in[18]
  PIN pc_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 796.000 694.970 800.000 ;
    END
  END pc_in[19]
  PIN pc_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END pc_in[1]
  PIN pc_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 796.000 600.210 800.000 ;
    END
  END pc_in[20]
  PIN pc_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 796.000 772.250 800.000 ;
    END
  END pc_in[21]
  PIN pc_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 796.000 487.970 800.000 ;
    END
  END pc_in[22]
  PIN pc_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 796.000 18.770 800.000 ;
    END
  END pc_in[23]
  PIN pc_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 796.000 746.490 800.000 ;
    END
  END pc_in[24]
  PIN pc_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 796.000 738.210 800.000 ;
    END
  END pc_in[25]
  PIN pc_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END pc_in[26]
  PIN pc_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END pc_in[27]
  PIN pc_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END pc_in[28]
  PIN pc_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END pc_in[29]
  PIN pc_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END pc_in[2]
  PIN pc_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 0.000 675.650 4.000 ;
    END
  END pc_in[30]
  PIN pc_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 796.000 105.250 800.000 ;
    END
  END pc_in[31]
  PIN pc_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END pc_in[3]
  PIN pc_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END pc_in[4]
  PIN pc_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 796.000 785.130 800.000 ;
    END
  END pc_in[5]
  PIN pc_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END pc_in[6]
  PIN pc_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 108.840 800.000 109.440 ;
    END
  END pc_in[7]
  PIN pc_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 796.000 96.050 800.000 ;
    END
  END pc_in[8]
  PIN pc_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 796.000 147.570 800.000 ;
    END
  END pc_in[9]
  PIN pc_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END pc_out[0]
  PIN pc_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 140.120 800.000 140.720 ;
    END
  END pc_out[10]
  PIN pc_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 796.000 126.410 800.000 ;
    END
  END pc_out[11]
  PIN pc_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 776.600 800.000 777.200 ;
    END
  END pc_out[12]
  PIN pc_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 63.960 800.000 64.560 ;
    END
  END pc_out[13]
  PIN pc_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END pc_out[14]
  PIN pc_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END pc_out[15]
  PIN pc_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 451.560 800.000 452.160 ;
    END
  END pc_out[16]
  PIN pc_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END pc_out[17]
  PIN pc_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 738.520 800.000 739.120 ;
    END
  END pc_out[18]
  PIN pc_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 572.600 800.000 573.200 ;
    END
  END pc_out[19]
  PIN pc_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END pc_out[1]
  PIN pc_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END pc_out[20]
  PIN pc_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 796.000 349.970 800.000 ;
    END
  END pc_out[21]
  PIN pc_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END pc_out[22]
  PIN pc_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 796.000 431.850 800.000 ;
    END
  END pc_out[23]
  PIN pc_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 70.760 800.000 71.360 ;
    END
  END pc_out[24]
  PIN pc_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END pc_out[25]
  PIN pc_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END pc_out[26]
  PIN pc_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END pc_out[27]
  PIN pc_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 796.000 492.570 800.000 ;
    END
  END pc_out[28]
  PIN pc_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 382.200 800.000 382.800 ;
    END
  END pc_out[29]
  PIN pc_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END pc_out[2]
  PIN pc_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 273.400 800.000 274.000 ;
    END
  END pc_out[30]
  PIN pc_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 4.000 ;
    END
  END pc_out[31]
  PIN pc_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END pc_out[3]
  PIN pc_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 267.960 800.000 268.560 ;
    END
  END pc_out[4]
  PIN pc_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END pc_out[5]
  PIN pc_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 12.280 800.000 12.880 ;
    END
  END pc_out[6]
  PIN pc_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END pc_out[7]
  PIN pc_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 76.200 800.000 76.800 ;
    END
  END pc_out[8]
  PIN pc_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 796.000 587.330 800.000 ;
    END
  END pc_out[9]
  PIN psw_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END psw_in
  PIN read_interactive_value_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 796.000 518.330 800.000 ;
    END
  END read_interactive_value_in[0]
  PIN read_interactive_value_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 796.000 638.850 800.000 ;
    END
  END read_interactive_value_in[10]
  PIN read_interactive_value_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END read_interactive_value_in[11]
  PIN read_interactive_value_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 796.000 118.130 800.000 ;
    END
  END read_interactive_value_in[12]
  PIN read_interactive_value_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 796.000 134.690 800.000 ;
    END
  END read_interactive_value_in[13]
  PIN read_interactive_value_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END read_interactive_value_in[14]
  PIN read_interactive_value_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END read_interactive_value_in[15]
  PIN read_interactive_value_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 432.520 800.000 433.120 ;
    END
  END read_interactive_value_in[16]
  PIN read_interactive_value_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END read_interactive_value_in[17]
  PIN read_interactive_value_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 413.480 800.000 414.080 ;
    END
  END read_interactive_value_in[18]
  PIN read_interactive_value_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END read_interactive_value_in[19]
  PIN read_interactive_value_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 796.000 229.450 800.000 ;
    END
  END read_interactive_value_in[1]
  PIN read_interactive_value_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 185.000 800.000 185.600 ;
    END
  END read_interactive_value_in[20]
  PIN read_interactive_value_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END read_interactive_value_in[21]
  PIN read_interactive_value_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 191.800 800.000 192.400 ;
    END
  END read_interactive_value_in[22]
  PIN read_interactive_value_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END read_interactive_value_in[23]
  PIN read_interactive_value_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 796.000 479.690 800.000 ;
    END
  END read_interactive_value_in[24]
  PIN read_interactive_value_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 363.160 800.000 363.760 ;
    END
  END read_interactive_value_in[25]
  PIN read_interactive_value_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END read_interactive_value_in[26]
  PIN read_interactive_value_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 796.000 418.970 800.000 ;
    END
  END read_interactive_value_in[27]
  PIN read_interactive_value_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END read_interactive_value_in[28]
  PIN read_interactive_value_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END read_interactive_value_in[29]
  PIN read_interactive_value_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 796.000 333.410 800.000 ;
    END
  END read_interactive_value_in[2]
  PIN read_interactive_value_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 629.720 800.000 630.320 ;
    END
  END read_interactive_value_in[30]
  PIN read_interactive_value_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 121.080 800.000 121.680 ;
    END
  END read_interactive_value_in[31]
  PIN read_interactive_value_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 669.160 800.000 669.760 ;
    END
  END read_interactive_value_in[3]
  PIN read_interactive_value_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END read_interactive_value_in[4]
  PIN read_interactive_value_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END read_interactive_value_in[5]
  PIN read_interactive_value_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END read_interactive_value_in[6]
  PIN read_interactive_value_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 489.640 800.000 490.240 ;
    END
  END read_interactive_value_in[7]
  PIN read_interactive_value_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 579.400 800.000 580.000 ;
    END
  END read_interactive_value_in[8]
  PIN read_interactive_value_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 796.000 14.170 800.000 ;
    END
  END read_interactive_value_in[9]
  PIN read_interactive_value_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END read_interactive_value_out[0]
  PIN read_interactive_value_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END read_interactive_value_out[10]
  PIN read_interactive_value_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 796.000 177.930 800.000 ;
    END
  END read_interactive_value_out[11]
  PIN read_interactive_value_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 38.120 800.000 38.720 ;
    END
  END read_interactive_value_out[12]
  PIN read_interactive_value_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END read_interactive_value_out[13]
  PIN read_interactive_value_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 796.000 457.610 800.000 ;
    END
  END read_interactive_value_out[14]
  PIN read_interactive_value_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.760 4.000 751.360 ;
    END
  END read_interactive_value_out[15]
  PIN read_interactive_value_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 750.760 800.000 751.360 ;
    END
  END read_interactive_value_out[16]
  PIN read_interactive_value_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 796.000 444.730 800.000 ;
    END
  END read_interactive_value_out[17]
  PIN read_interactive_value_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END read_interactive_value_out[18]
  PIN read_interactive_value_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END read_interactive_value_out[19]
  PIN read_interactive_value_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END read_interactive_value_out[1]
  PIN read_interactive_value_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END read_interactive_value_out[20]
  PIN read_interactive_value_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 439.320 800.000 439.920 ;
    END
  END read_interactive_value_out[21]
  PIN read_interactive_value_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 796.000 303.050 800.000 ;
    END
  END read_interactive_value_out[22]
  PIN read_interactive_value_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 688.200 800.000 688.800 ;
    END
  END read_interactive_value_out[23]
  PIN read_interactive_value_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 796.000 5.890 800.000 ;
    END
  END read_interactive_value_out[24]
  PIN read_interactive_value_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 796.000 604.810 800.000 ;
    END
  END read_interactive_value_out[25]
  PIN read_interactive_value_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 605.240 800.000 605.840 ;
    END
  END read_interactive_value_out[26]
  PIN read_interactive_value_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 796.000 290.170 800.000 ;
    END
  END read_interactive_value_out[27]
  PIN read_interactive_value_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 731.720 800.000 732.320 ;
    END
  END read_interactive_value_out[28]
  PIN read_interactive_value_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 796.000 337.090 800.000 ;
    END
  END read_interactive_value_out[29]
  PIN read_interactive_value_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END read_interactive_value_out[2]
  PIN read_interactive_value_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END read_interactive_value_out[30]
  PIN read_interactive_value_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 31.320 800.000 31.920 ;
    END
  END read_interactive_value_out[31]
  PIN read_interactive_value_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END read_interactive_value_out[3]
  PIN read_interactive_value_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 796.000 556.970 800.000 ;
    END
  END read_interactive_value_out[4]
  PIN read_interactive_value_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 796.000 643.450 800.000 ;
    END
  END read_interactive_value_out[5]
  PIN read_interactive_value_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END read_interactive_value_out[6]
  PIN read_interactive_value_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 89.800 800.000 90.400 ;
    END
  END read_interactive_value_out[7]
  PIN read_interactive_value_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 796.000 143.890 800.000 ;
    END
  END read_interactive_value_out[8]
  PIN read_interactive_value_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 796.000 195.410 800.000 ;
    END
  END read_interactive_value_out[9]
  PIN reg_data_alu_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 796.000 393.210 800.000 ;
    END
  END reg_data_alu_in[0]
  PIN reg_data_alu_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END reg_data_alu_in[10]
  PIN reg_data_alu_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 796.000 428.170 800.000 ;
    END
  END reg_data_alu_in[11]
  PIN reg_data_alu_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 306.040 800.000 306.640 ;
    END
  END reg_data_alu_in[12]
  PIN reg_data_alu_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END reg_data_alu_in[13]
  PIN reg_data_alu_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END reg_data_alu_in[14]
  PIN reg_data_alu_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 796.000 113.530 800.000 ;
    END
  END reg_data_alu_in[15]
  PIN reg_data_alu_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END reg_data_alu_in[16]
  PIN reg_data_alu_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 19.080 800.000 19.680 ;
    END
  END reg_data_alu_in[17]
  PIN reg_data_alu_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 693.640 800.000 694.240 ;
    END
  END reg_data_alu_in[18]
  PIN reg_data_alu_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END reg_data_alu_in[19]
  PIN reg_data_alu_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END reg_data_alu_in[1]
  PIN reg_data_alu_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 796.000 751.090 800.000 ;
    END
  END reg_data_alu_in[20]
  PIN reg_data_alu_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 369.960 800.000 370.560 ;
    END
  END reg_data_alu_in[21]
  PIN reg_data_alu_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 229.880 800.000 230.480 ;
    END
  END reg_data_alu_in[22]
  PIN reg_data_alu_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END reg_data_alu_in[23]
  PIN reg_data_alu_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 796.000 92.370 800.000 ;
    END
  END reg_data_alu_in[24]
  PIN reg_data_alu_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END reg_data_alu_in[25]
  PIN reg_data_alu_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 796.000 346.290 800.000 ;
    END
  END reg_data_alu_in[26]
  PIN reg_data_alu_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END reg_data_alu_in[27]
  PIN reg_data_alu_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END reg_data_alu_in[28]
  PIN reg_data_alu_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END reg_data_alu_in[29]
  PIN reg_data_alu_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END reg_data_alu_in[2]
  PIN reg_data_alu_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END reg_data_alu_in[30]
  PIN reg_data_alu_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 788.840 800.000 789.440 ;
    END
  END reg_data_alu_in[31]
  PIN reg_data_alu_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 796.000 187.130 800.000 ;
    END
  END reg_data_alu_in[3]
  PIN reg_data_alu_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END reg_data_alu_in[4]
  PIN reg_data_alu_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 796.000 685.770 800.000 ;
    END
  END reg_data_alu_in[5]
  PIN reg_data_alu_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 796.000 500.850 800.000 ;
    END
  END reg_data_alu_in[6]
  PIN reg_data_alu_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 197.240 800.000 197.840 ;
    END
  END reg_data_alu_in[7]
  PIN reg_data_alu_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END reg_data_alu_in[8]
  PIN reg_data_alu_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 796.000 62.010 800.000 ;
    END
  END reg_data_alu_in[9]
  PIN reg_data_alu_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 681.400 800.000 682.000 ;
    END
  END reg_data_alu_out[0]
  PIN reg_data_alu_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 796.000 131.010 800.000 ;
    END
  END reg_data_alu_out[10]
  PIN reg_data_alu_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END reg_data_alu_out[11]
  PIN reg_data_alu_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 796.000 307.650 800.000 ;
    END
  END reg_data_alu_out[12]
  PIN reg_data_alu_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END reg_data_alu_out[13]
  PIN reg_data_alu_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END reg_data_alu_out[14]
  PIN reg_data_alu_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END reg_data_alu_out[15]
  PIN reg_data_alu_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 796.000 754.770 800.000 ;
    END
  END reg_data_alu_out[16]
  PIN reg_data_alu_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 95.240 800.000 95.840 ;
    END
  END reg_data_alu_out[17]
  PIN reg_data_alu_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END reg_data_alu_out[18]
  PIN reg_data_alu_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END reg_data_alu_out[19]
  PIN reg_data_alu_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 796.000 255.210 800.000 ;
    END
  END reg_data_alu_out[1]
  PIN reg_data_alu_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 796.000 74.890 800.000 ;
    END
  END reg_data_alu_out[20]
  PIN reg_data_alu_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END reg_data_alu_out[21]
  PIN reg_data_alu_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END reg_data_alu_out[22]
  PIN reg_data_alu_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 344.120 800.000 344.720 ;
    END
  END reg_data_alu_out[23]
  PIN reg_data_alu_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 796.000 375.730 800.000 ;
    END
  END reg_data_alu_out[24]
  PIN reg_data_alu_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 318.280 800.000 318.880 ;
    END
  END reg_data_alu_out[25]
  PIN reg_data_alu_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END reg_data_alu_out[26]
  PIN reg_data_alu_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END reg_data_alu_out[27]
  PIN reg_data_alu_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END reg_data_alu_out[28]
  PIN reg_data_alu_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END reg_data_alu_out[29]
  PIN reg_data_alu_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 796.000 272.690 800.000 ;
    END
  END reg_data_alu_out[2]
  PIN reg_data_alu_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END reg_data_alu_out[30]
  PIN reg_data_alu_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END reg_data_alu_out[31]
  PIN reg_data_alu_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 796.000 79.490 800.000 ;
    END
  END reg_data_alu_out[3]
  PIN reg_data_alu_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 796.000 264.410 800.000 ;
    END
  END reg_data_alu_out[4]
  PIN reg_data_alu_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END reg_data_alu_out[5]
  PIN reg_data_alu_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END reg_data_alu_out[6]
  PIN reg_data_alu_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END reg_data_alu_out[7]
  PIN reg_data_alu_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END reg_data_alu_out[8]
  PIN reg_data_alu_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END reg_data_alu_out[9]
  PIN reg_dest_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 796.000 703.250 800.000 ;
    END
  END reg_dest_in[0]
  PIN reg_dest_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END reg_dest_in[1]
  PIN reg_dest_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 796.000 328.810 800.000 ;
    END
  END reg_dest_in[2]
  PIN reg_dest_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END reg_dest_in[3]
  PIN reg_dest_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 796.000 173.330 800.000 ;
    END
  END reg_dest_in[4]
  PIN reg_dest_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 796.000 372.050 800.000 ;
    END
  END reg_dest_out[0]
  PIN reg_dest_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END reg_dest_out[1]
  PIN reg_dest_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END reg_dest_out[2]
  PIN reg_dest_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 796.000 169.650 800.000 ;
    END
  END reg_dest_out[3]
  PIN reg_dest_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 51.720 800.000 52.320 ;
    END
  END reg_dest_out[4]
  PIN reg_write_enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 0.040 800.000 0.640 ;
    END
  END reg_write_enable_in
  PIN reg_write_enable_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END reg_write_enable_out
  PIN rm0_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 796.000 57.410 800.000 ;
    END
  END rm0_in[0]
  PIN rm0_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END rm0_in[10]
  PIN rm0_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 796.000 776.850 800.000 ;
    END
  END rm0_in[11]
  PIN rm0_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END rm0_in[12]
  PIN rm0_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END rm0_in[13]
  PIN rm0_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END rm0_in[14]
  PIN rm0_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 4.000 ;
    END
  END rm0_in[15]
  PIN rm0_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 356.360 800.000 356.960 ;
    END
  END rm0_in[16]
  PIN rm0_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 796.000 466.810 800.000 ;
    END
  END rm0_in[17]
  PIN rm0_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 796.000 367.450 800.000 ;
    END
  END rm0_in[18]
  PIN rm0_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END rm0_in[19]
  PIN rm0_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 796.000 156.770 800.000 ;
    END
  END rm0_in[1]
  PIN rm0_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END rm0_in[20]
  PIN rm0_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 796.000 27.050 800.000 ;
    END
  END rm0_in[21]
  PIN rm0_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 796.000 672.890 800.000 ;
    END
  END rm0_in[22]
  PIN rm0_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END rm0_in[23]
  PIN rm0_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 796.000 384.930 800.000 ;
    END
  END rm0_in[24]
  PIN rm0_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END rm0_in[25]
  PIN rm0_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 133.320 800.000 133.920 ;
    END
  END rm0_in[26]
  PIN rm0_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 796.000 677.490 800.000 ;
    END
  END rm0_in[27]
  PIN rm0_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 796.000 656.330 800.000 ;
    END
  END rm0_in[28]
  PIN rm0_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END rm0_in[29]
  PIN rm0_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END rm0_in[2]
  PIN rm0_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 796.000 320.530 800.000 ;
    END
  END rm0_in[30]
  PIN rm0_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 796.000 246.930 800.000 ;
    END
  END rm0_in[31]
  PIN rm0_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END rm0_in[3]
  PIN rm0_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END rm0_in[4]
  PIN rm0_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END rm0_in[5]
  PIN rm0_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 796.000 225.770 800.000 ;
    END
  END rm0_in[6]
  PIN rm0_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END rm0_in[7]
  PIN rm0_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 796.000 763.970 800.000 ;
    END
  END rm0_in[8]
  PIN rm0_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 394.440 800.000 395.040 ;
    END
  END rm0_in[9]
  PIN rm0_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 796.000 548.690 800.000 ;
    END
  END rm0_out[0]
  PIN rm0_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 796.000 625.970 800.000 ;
    END
  END rm0_out[10]
  PIN rm0_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END rm0_out[11]
  PIN rm0_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 591.640 800.000 592.240 ;
    END
  END rm0_out[12]
  PIN rm0_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 4.000 ;
    END
  END rm0_out[13]
  PIN rm0_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 350.920 800.000 351.520 ;
    END
  END rm0_out[14]
  PIN rm0_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END rm0_out[15]
  PIN rm0_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END rm0_out[16]
  PIN rm0_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END rm0_out[17]
  PIN rm0_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END rm0_out[18]
  PIN rm0_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END rm0_out[19]
  PIN rm0_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 223.080 800.000 223.680 ;
    END
  END rm0_out[1]
  PIN rm0_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END rm0_out[20]
  PIN rm0_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 401.240 800.000 401.840 ;
    END
  END rm0_out[21]
  PIN rm0_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 796.000 268.090 800.000 ;
    END
  END rm0_out[22]
  PIN rm0_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END rm0_out[23]
  PIN rm0_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 796.000 522.930 800.000 ;
    END
  END rm0_out[24]
  PIN rm0_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 655.560 800.000 656.160 ;
    END
  END rm0_out[25]
  PIN rm0_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END rm0_out[26]
  PIN rm0_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 311.480 800.000 312.080 ;
    END
  END rm0_out[27]
  PIN rm0_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END rm0_out[28]
  PIN rm0_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 83.000 800.000 83.600 ;
    END
  END rm0_out[29]
  PIN rm0_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 796.000 23.370 800.000 ;
    END
  END rm0_out[2]
  PIN rm0_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 796.000 513.730 800.000 ;
    END
  END rm0_out[30]
  PIN rm0_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END rm0_out[31]
  PIN rm0_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END rm0_out[3]
  PIN rm0_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.120 4.000 718.720 ;
    END
  END rm0_out[4]
  PIN rm0_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 6.840 800.000 7.440 ;
    END
  END rm0_out[5]
  PIN rm0_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END rm0_out[6]
  PIN rm0_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END rm0_out[7]
  PIN rm0_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 4.000 ;
    END
  END rm0_out[8]
  PIN rm0_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 757.560 800.000 758.160 ;
    END
  END rm0_out[9]
  PIN rm1_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END rm1_in[0]
  PIN rm1_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END rm1_in[10]
  PIN rm1_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 171.400 800.000 172.000 ;
    END
  END rm1_in[11]
  PIN rm1_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END rm1_in[12]
  PIN rm1_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 796.000 100.650 800.000 ;
    END
  END rm1_in[13]
  PIN rm1_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END rm1_in[14]
  PIN rm1_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 375.400 800.000 376.000 ;
    END
  END rm1_in[15]
  PIN rm1_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 796.000 780.530 800.000 ;
    END
  END rm1_in[16]
  PIN rm1_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 796.000 707.850 800.000 ;
    END
  END rm1_in[17]
  PIN rm1_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END rm1_in[18]
  PIN rm1_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 796.000 789.730 800.000 ;
    END
  END rm1_in[19]
  PIN rm1_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 796.000 294.770 800.000 ;
    END
  END rm1_in[1]
  PIN rm1_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END rm1_in[20]
  PIN rm1_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END rm1_in[21]
  PIN rm1_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 152.360 800.000 152.960 ;
    END
  END rm1_in[22]
  PIN rm1_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 408.040 800.000 408.640 ;
    END
  END rm1_in[23]
  PIN rm1_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 796.000 436.450 800.000 ;
    END
  END rm1_in[24]
  PIN rm1_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END rm1_in[25]
  PIN rm1_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 636.520 800.000 637.120 ;
    END
  END rm1_in[26]
  PIN rm1_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 510.040 800.000 510.640 ;
    END
  END rm1_in[27]
  PIN rm1_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 796.000 725.330 800.000 ;
    END
  END rm1_in[28]
  PIN rm1_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 726.280 800.000 726.880 ;
    END
  END rm1_in[29]
  PIN rm1_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END rm1_in[2]
  PIN rm1_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 796.000 139.290 800.000 ;
    END
  END rm1_in[30]
  PIN rm1_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END rm1_in[31]
  PIN rm1_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END rm1_in[3]
  PIN rm1_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END rm1_in[4]
  PIN rm1_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END rm1_in[5]
  PIN rm1_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END rm1_in[6]
  PIN rm1_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 127.880 800.000 128.480 ;
    END
  END rm1_in[7]
  PIN rm1_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 643.320 800.000 643.920 ;
    END
  END rm1_in[8]
  PIN rm1_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END rm1_in[9]
  PIN rm1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 796.000 423.570 800.000 ;
    END
  END rm1_out[0]
  PIN rm1_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 796.000 315.930 800.000 ;
    END
  END rm1_out[10]
  PIN rm1_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END rm1_out[11]
  PIN rm1_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 745.320 800.000 745.920 ;
    END
  END rm1_out[12]
  PIN rm1_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END rm1_out[13]
  PIN rm1_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END rm1_out[14]
  PIN rm1_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END rm1_out[15]
  PIN rm1_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 624.280 800.000 624.880 ;
    END
  END rm1_out[16]
  PIN rm1_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 796.000 578.130 800.000 ;
    END
  END rm1_out[17]
  PIN rm1_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 796.000 65.690 800.000 ;
    END
  END rm1_out[18]
  PIN rm1_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 796.000 660.010 800.000 ;
    END
  END rm1_out[19]
  PIN rm1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 796.000 690.370 800.000 ;
    END
  END rm1_out[1]
  PIN rm1_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END rm1_out[20]
  PIN rm1_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END rm1_out[21]
  PIN rm1_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 796.000 470.490 800.000 ;
    END
  END rm1_out[22]
  PIN rm1_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END rm1_out[23]
  PIN rm1_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END rm1_out[24]
  PIN rm1_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END rm1_out[25]
  PIN rm1_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END rm1_out[26]
  PIN rm1_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 25.880 800.000 26.480 ;
    END
  END rm1_out[27]
  PIN rm1_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 796.000 539.490 800.000 ;
    END
  END rm1_out[28]
  PIN rm1_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END rm1_out[29]
  PIN rm1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END rm1_out[2]
  PIN rm1_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END rm1_out[30]
  PIN rm1_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END rm1_out[31]
  PIN rm1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END rm1_out[3]
  PIN rm1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 796.000 453.930 800.000 ;
    END
  END rm1_out[4]
  PIN rm1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END rm1_out[5]
  PIN rm1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END rm1_out[6]
  PIN rm1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END rm1_out[7]
  PIN rm1_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END rm1_out[8]
  PIN rm1_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 719.480 800.000 720.080 ;
    END
  END rm1_out[9]
  PIN rm2_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END rm2_in[0]
  PIN rm2_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END rm2_in[10]
  PIN rm2_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 0.000 762.130 4.000 ;
    END
  END rm2_in[11]
  PIN rm2_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END rm2_in[12]
  PIN rm2_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 796.000 362.850 800.000 ;
    END
  END rm2_in[13]
  PIN rm2_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 529.080 800.000 529.680 ;
    END
  END rm2_in[14]
  PIN rm2_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END rm2_in[15]
  PIN rm2_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 796.000 526.610 800.000 ;
    END
  END rm2_in[16]
  PIN rm2_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 57.160 800.000 57.760 ;
    END
  END rm2_in[17]
  PIN rm2_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 796.000 311.330 800.000 ;
    END
  END rm2_in[18]
  PIN rm2_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END rm2_in[19]
  PIN rm2_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 796.000 49.130 800.000 ;
    END
  END rm2_in[1]
  PIN rm2_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END rm2_in[20]
  PIN rm2_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END rm2_in[21]
  PIN rm2_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END rm2_in[22]
  PIN rm2_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 662.360 800.000 662.960 ;
    END
  END rm2_in[23]
  PIN rm2_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END rm2_in[24]
  PIN rm2_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END rm2_in[25]
  PIN rm2_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 796.000 108.930 800.000 ;
    END
  END rm2_in[26]
  PIN rm2_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 796.000 535.810 800.000 ;
    END
  END rm2_in[27]
  PIN rm2_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 769.800 800.000 770.400 ;
    END
  END rm2_in[28]
  PIN rm2_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 796.000 83.170 800.000 ;
    END
  END rm2_in[29]
  PIN rm2_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 796.000 152.170 800.000 ;
    END
  END rm2_in[2]
  PIN rm2_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 114.280 800.000 114.880 ;
    END
  END rm2_in[30]
  PIN rm2_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 796.000 44.530 800.000 ;
    END
  END rm2_in[31]
  PIN rm2_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END rm2_in[3]
  PIN rm2_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 796.000 406.090 800.000 ;
    END
  END rm2_in[4]
  PIN rm2_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 796.000 251.530 800.000 ;
    END
  END rm2_in[5]
  PIN rm2_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END rm2_in[6]
  PIN rm2_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END rm2_in[7]
  PIN rm2_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END rm2_in[8]
  PIN rm2_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 712.680 800.000 713.280 ;
    END
  END rm2_in[9]
  PIN rm2_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 650.120 800.000 650.720 ;
    END
  END rm2_out[0]
  PIN rm2_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END rm2_out[10]
  PIN rm2_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 567.160 800.000 567.760 ;
    END
  END rm2_out[11]
  PIN rm2_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 248.920 800.000 249.520 ;
    END
  END rm2_out[12]
  PIN rm2_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END rm2_out[13]
  PIN rm2_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 796.000 415.290 800.000 ;
    END
  END rm2_out[14]
  PIN rm2_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END rm2_out[15]
  PIN rm2_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END rm2_out[16]
  PIN rm2_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END rm2_out[17]
  PIN rm2_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 146.920 800.000 147.520 ;
    END
  END rm2_out[18]
  PIN rm2_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 796.000 39.930 800.000 ;
    END
  END rm2_out[19]
  PIN rm2_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END rm2_out[1]
  PIN rm2_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END rm2_out[20]
  PIN rm2_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END rm2_out[21]
  PIN rm2_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 515.480 800.000 516.080 ;
    END
  END rm2_out[22]
  PIN rm2_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 796.000 720.730 800.000 ;
    END
  END rm2_out[23]
  PIN rm2_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END rm2_out[24]
  PIN rm2_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 796.000 544.090 800.000 ;
    END
  END rm2_out[25]
  PIN rm2_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 337.320 800.000 337.920 ;
    END
  END rm2_out[26]
  PIN rm2_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END rm2_out[27]
  PIN rm2_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 796.000 531.210 800.000 ;
    END
  END rm2_out[28]
  PIN rm2_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END rm2_out[29]
  PIN rm2_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END rm2_out[2]
  PIN rm2_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END rm2_out[30]
  PIN rm2_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END rm2_out[31]
  PIN rm2_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 165.960 800.000 166.560 ;
    END
  END rm2_out[3]
  PIN rm2_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 796.000 216.570 800.000 ;
    END
  END rm2_out[4]
  PIN rm2_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 796.000 798.010 800.000 ;
    END
  END rm2_out[5]
  PIN rm2_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END rm2_out[6]
  PIN rm2_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END rm2_out[7]
  PIN rm2_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END rm2_out[8]
  PIN rm2_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END rm2_out[9]
  PIN stall
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END stall
  PIN stored_rm4_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 420.280 800.000 420.880 ;
    END
  END stored_rm4_in[0]
  PIN stored_rm4_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END stored_rm4_in[10]
  PIN stored_rm4_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 796.000 497.170 800.000 ;
    END
  END stored_rm4_in[11]
  PIN stored_rm4_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 796.000 669.210 800.000 ;
    END
  END stored_rm4_in[12]
  PIN stored_rm4_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 796.000 52.810 800.000 ;
    END
  END stored_rm4_in[13]
  PIN stored_rm4_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END stored_rm4_in[14]
  PIN stored_rm4_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 496.440 800.000 497.040 ;
    END
  END stored_rm4_in[15]
  PIN stored_rm4_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 796.000 699.570 800.000 ;
    END
  END stored_rm4_in[16]
  PIN stored_rm4_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END stored_rm4_in[17]
  PIN stored_rm4_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 674.600 800.000 675.200 ;
    END
  END stored_rm4_in[18]
  PIN stored_rm4_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 204.040 800.000 204.640 ;
    END
  END stored_rm4_in[19]
  PIN stored_rm4_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END stored_rm4_in[1]
  PIN stored_rm4_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 796.000 621.370 800.000 ;
    END
  END stored_rm4_in[20]
  PIN stored_rm4_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 796.000 208.290 800.000 ;
    END
  END stored_rm4_in[21]
  PIN stored_rm4_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END stored_rm4_in[22]
  PIN stored_rm4_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 484.200 800.000 484.800 ;
    END
  END stored_rm4_in[23]
  PIN stored_rm4_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END stored_rm4_in[24]
  PIN stored_rm4_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 159.160 800.000 159.760 ;
    END
  END stored_rm4_in[25]
  PIN stored_rm4_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END stored_rm4_in[26]
  PIN stored_rm4_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END stored_rm4_in[27]
  PIN stored_rm4_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END stored_rm4_in[28]
  PIN stored_rm4_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END stored_rm4_in[29]
  PIN stored_rm4_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 292.440 800.000 293.040 ;
    END
  END stored_rm4_in[2]
  PIN stored_rm4_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 796.000 608.490 800.000 ;
    END
  END stored_rm4_in[30]
  PIN stored_rm4_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 764.360 800.000 764.960 ;
    END
  END stored_rm4_in[31]
  PIN stored_rm4_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END stored_rm4_in[3]
  PIN stored_rm4_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END stored_rm4_in[4]
  PIN stored_rm4_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 427.080 800.000 427.680 ;
    END
  END stored_rm4_in[5]
  PIN stored_rm4_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END stored_rm4_in[6]
  PIN stored_rm4_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 783.400 800.000 784.000 ;
    END
  END stored_rm4_in[7]
  PIN stored_rm4_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 796.000 591.010 800.000 ;
    END
  END stored_rm4_in[8]
  PIN stored_rm4_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END stored_rm4_in[9]
  PIN stored_rm4_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 796.000 569.850 800.000 ;
    END
  END stored_rm4_out[0]
  PIN stored_rm4_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END stored_rm4_out[10]
  PIN stored_rm4_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END stored_rm4_out[11]
  PIN stored_rm4_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END stored_rm4_out[12]
  PIN stored_rm4_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END stored_rm4_out[13]
  PIN stored_rm4_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 0.000 542.250 4.000 ;
    END
  END stored_rm4_out[14]
  PIN stored_rm4_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END stored_rm4_out[15]
  PIN stored_rm4_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END stored_rm4_out[16]
  PIN stored_rm4_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 796.000 277.290 800.000 ;
    END
  END stored_rm4_out[17]
  PIN stored_rm4_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END stored_rm4_out[18]
  PIN stored_rm4_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END stored_rm4_out[19]
  PIN stored_rm4_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END stored_rm4_out[1]
  PIN stored_rm4_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 796.000 449.330 800.000 ;
    END
  END stored_rm4_out[20]
  PIN stored_rm4_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 796.000 298.450 800.000 ;
    END
  END stored_rm4_out[21]
  PIN stored_rm4_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END stored_rm4_out[22]
  PIN stored_rm4_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 796.000 574.450 800.000 ;
    END
  END stored_rm4_out[23]
  PIN stored_rm4_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 102.040 800.000 102.640 ;
    END
  END stored_rm4_out[24]
  PIN stored_rm4_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END stored_rm4_out[25]
  PIN stored_rm4_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 598.440 800.000 599.040 ;
    END
  END stored_rm4_out[26]
  PIN stored_rm4_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END stored_rm4_out[27]
  PIN stored_rm4_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END stored_rm4_out[28]
  PIN stored_rm4_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END stored_rm4_out[29]
  PIN stored_rm4_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 553.560 800.000 554.160 ;
    END
  END stored_rm4_out[2]
  PIN stored_rm4_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END stored_rm4_out[30]
  PIN stored_rm4_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 796.000 561.570 800.000 ;
    END
  END stored_rm4_out[31]
  PIN stored_rm4_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 796.000 552.370 800.000 ;
    END
  END stored_rm4_out[3]
  PIN stored_rm4_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 796.000 70.290 800.000 ;
    END
  END stored_rm4_out[4]
  PIN stored_rm4_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 796.000 190.810 800.000 ;
    END
  END stored_rm4_out[5]
  PIN stored_rm4_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END stored_rm4_out[6]
  PIN stored_rm4_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END stored_rm4_out[7]
  PIN stored_rm4_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 796.000 10.490 800.000 ;
    END
  END stored_rm4_out[8]
  PIN stored_rm4_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 299.240 800.000 299.840 ;
    END
  END stored_rm4_out[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 0.425 797.035 795.855 ;
      LAYER met1 ;
        RECT 0.070 0.380 798.030 795.900 ;
      LAYER met2 ;
        RECT 0.100 795.720 0.730 796.690 ;
        RECT 1.570 795.720 5.330 796.690 ;
        RECT 6.170 795.720 9.930 796.690 ;
        RECT 10.770 795.720 13.610 796.690 ;
        RECT 14.450 795.720 18.210 796.690 ;
        RECT 19.050 795.720 22.810 796.690 ;
        RECT 23.650 795.720 26.490 796.690 ;
        RECT 27.330 795.720 31.090 796.690 ;
        RECT 31.930 795.720 35.690 796.690 ;
        RECT 36.530 795.720 39.370 796.690 ;
        RECT 40.210 795.720 43.970 796.690 ;
        RECT 44.810 795.720 48.570 796.690 ;
        RECT 49.410 795.720 52.250 796.690 ;
        RECT 53.090 795.720 56.850 796.690 ;
        RECT 57.690 795.720 61.450 796.690 ;
        RECT 62.290 795.720 65.130 796.690 ;
        RECT 65.970 795.720 69.730 796.690 ;
        RECT 70.570 795.720 74.330 796.690 ;
        RECT 75.170 795.720 78.930 796.690 ;
        RECT 79.770 795.720 82.610 796.690 ;
        RECT 83.450 795.720 87.210 796.690 ;
        RECT 88.050 795.720 91.810 796.690 ;
        RECT 92.650 795.720 95.490 796.690 ;
        RECT 96.330 795.720 100.090 796.690 ;
        RECT 100.930 795.720 104.690 796.690 ;
        RECT 105.530 795.720 108.370 796.690 ;
        RECT 109.210 795.720 112.970 796.690 ;
        RECT 113.810 795.720 117.570 796.690 ;
        RECT 118.410 795.720 121.250 796.690 ;
        RECT 122.090 795.720 125.850 796.690 ;
        RECT 126.690 795.720 130.450 796.690 ;
        RECT 131.290 795.720 134.130 796.690 ;
        RECT 134.970 795.720 138.730 796.690 ;
        RECT 139.570 795.720 143.330 796.690 ;
        RECT 144.170 795.720 147.010 796.690 ;
        RECT 147.850 795.720 151.610 796.690 ;
        RECT 152.450 795.720 156.210 796.690 ;
        RECT 157.050 795.720 159.890 796.690 ;
        RECT 160.730 795.720 164.490 796.690 ;
        RECT 165.330 795.720 169.090 796.690 ;
        RECT 169.930 795.720 172.770 796.690 ;
        RECT 173.610 795.720 177.370 796.690 ;
        RECT 178.210 795.720 181.970 796.690 ;
        RECT 182.810 795.720 186.570 796.690 ;
        RECT 187.410 795.720 190.250 796.690 ;
        RECT 191.090 795.720 194.850 796.690 ;
        RECT 195.690 795.720 199.450 796.690 ;
        RECT 200.290 795.720 203.130 796.690 ;
        RECT 203.970 795.720 207.730 796.690 ;
        RECT 208.570 795.720 212.330 796.690 ;
        RECT 213.170 795.720 216.010 796.690 ;
        RECT 216.850 795.720 220.610 796.690 ;
        RECT 221.450 795.720 225.210 796.690 ;
        RECT 226.050 795.720 228.890 796.690 ;
        RECT 229.730 795.720 233.490 796.690 ;
        RECT 234.330 795.720 238.090 796.690 ;
        RECT 238.930 795.720 241.770 796.690 ;
        RECT 242.610 795.720 246.370 796.690 ;
        RECT 247.210 795.720 250.970 796.690 ;
        RECT 251.810 795.720 254.650 796.690 ;
        RECT 255.490 795.720 259.250 796.690 ;
        RECT 260.090 795.720 263.850 796.690 ;
        RECT 264.690 795.720 267.530 796.690 ;
        RECT 268.370 795.720 272.130 796.690 ;
        RECT 272.970 795.720 276.730 796.690 ;
        RECT 277.570 795.720 280.410 796.690 ;
        RECT 281.250 795.720 285.010 796.690 ;
        RECT 285.850 795.720 289.610 796.690 ;
        RECT 290.450 795.720 294.210 796.690 ;
        RECT 295.050 795.720 297.890 796.690 ;
        RECT 298.730 795.720 302.490 796.690 ;
        RECT 303.330 795.720 307.090 796.690 ;
        RECT 307.930 795.720 310.770 796.690 ;
        RECT 311.610 795.720 315.370 796.690 ;
        RECT 316.210 795.720 319.970 796.690 ;
        RECT 320.810 795.720 323.650 796.690 ;
        RECT 324.490 795.720 328.250 796.690 ;
        RECT 329.090 795.720 332.850 796.690 ;
        RECT 333.690 795.720 336.530 796.690 ;
        RECT 337.370 795.720 341.130 796.690 ;
        RECT 341.970 795.720 345.730 796.690 ;
        RECT 346.570 795.720 349.410 796.690 ;
        RECT 350.250 795.720 354.010 796.690 ;
        RECT 354.850 795.720 358.610 796.690 ;
        RECT 359.450 795.720 362.290 796.690 ;
        RECT 363.130 795.720 366.890 796.690 ;
        RECT 367.730 795.720 371.490 796.690 ;
        RECT 372.330 795.720 375.170 796.690 ;
        RECT 376.010 795.720 379.770 796.690 ;
        RECT 380.610 795.720 384.370 796.690 ;
        RECT 385.210 795.720 388.970 796.690 ;
        RECT 389.810 795.720 392.650 796.690 ;
        RECT 393.490 795.720 397.250 796.690 ;
        RECT 398.090 795.720 401.850 796.690 ;
        RECT 402.690 795.720 405.530 796.690 ;
        RECT 406.370 795.720 410.130 796.690 ;
        RECT 410.970 795.720 414.730 796.690 ;
        RECT 415.570 795.720 418.410 796.690 ;
        RECT 419.250 795.720 423.010 796.690 ;
        RECT 423.850 795.720 427.610 796.690 ;
        RECT 428.450 795.720 431.290 796.690 ;
        RECT 432.130 795.720 435.890 796.690 ;
        RECT 436.730 795.720 440.490 796.690 ;
        RECT 441.330 795.720 444.170 796.690 ;
        RECT 445.010 795.720 448.770 796.690 ;
        RECT 449.610 795.720 453.370 796.690 ;
        RECT 454.210 795.720 457.050 796.690 ;
        RECT 457.890 795.720 461.650 796.690 ;
        RECT 462.490 795.720 466.250 796.690 ;
        RECT 467.090 795.720 469.930 796.690 ;
        RECT 470.770 795.720 474.530 796.690 ;
        RECT 475.370 795.720 479.130 796.690 ;
        RECT 479.970 795.720 482.810 796.690 ;
        RECT 483.650 795.720 487.410 796.690 ;
        RECT 488.250 795.720 492.010 796.690 ;
        RECT 492.850 795.720 496.610 796.690 ;
        RECT 497.450 795.720 500.290 796.690 ;
        RECT 501.130 795.720 504.890 796.690 ;
        RECT 505.730 795.720 509.490 796.690 ;
        RECT 510.330 795.720 513.170 796.690 ;
        RECT 514.010 795.720 517.770 796.690 ;
        RECT 518.610 795.720 522.370 796.690 ;
        RECT 523.210 795.720 526.050 796.690 ;
        RECT 526.890 795.720 530.650 796.690 ;
        RECT 531.490 795.720 535.250 796.690 ;
        RECT 536.090 795.720 538.930 796.690 ;
        RECT 539.770 795.720 543.530 796.690 ;
        RECT 544.370 795.720 548.130 796.690 ;
        RECT 548.970 795.720 551.810 796.690 ;
        RECT 552.650 795.720 556.410 796.690 ;
        RECT 557.250 795.720 561.010 796.690 ;
        RECT 561.850 795.720 564.690 796.690 ;
        RECT 565.530 795.720 569.290 796.690 ;
        RECT 570.130 795.720 573.890 796.690 ;
        RECT 574.730 795.720 577.570 796.690 ;
        RECT 578.410 795.720 582.170 796.690 ;
        RECT 583.010 795.720 586.770 796.690 ;
        RECT 587.610 795.720 590.450 796.690 ;
        RECT 591.290 795.720 595.050 796.690 ;
        RECT 595.890 795.720 599.650 796.690 ;
        RECT 600.490 795.720 604.250 796.690 ;
        RECT 605.090 795.720 607.930 796.690 ;
        RECT 608.770 795.720 612.530 796.690 ;
        RECT 613.370 795.720 617.130 796.690 ;
        RECT 617.970 795.720 620.810 796.690 ;
        RECT 621.650 795.720 625.410 796.690 ;
        RECT 626.250 795.720 630.010 796.690 ;
        RECT 630.850 795.720 633.690 796.690 ;
        RECT 634.530 795.720 638.290 796.690 ;
        RECT 639.130 795.720 642.890 796.690 ;
        RECT 643.730 795.720 646.570 796.690 ;
        RECT 647.410 795.720 651.170 796.690 ;
        RECT 652.010 795.720 655.770 796.690 ;
        RECT 656.610 795.720 659.450 796.690 ;
        RECT 660.290 795.720 664.050 796.690 ;
        RECT 664.890 795.720 668.650 796.690 ;
        RECT 669.490 795.720 672.330 796.690 ;
        RECT 673.170 795.720 676.930 796.690 ;
        RECT 677.770 795.720 681.530 796.690 ;
        RECT 682.370 795.720 685.210 796.690 ;
        RECT 686.050 795.720 689.810 796.690 ;
        RECT 690.650 795.720 694.410 796.690 ;
        RECT 695.250 795.720 699.010 796.690 ;
        RECT 699.850 795.720 702.690 796.690 ;
        RECT 703.530 795.720 707.290 796.690 ;
        RECT 708.130 795.720 711.890 796.690 ;
        RECT 712.730 795.720 715.570 796.690 ;
        RECT 716.410 795.720 720.170 796.690 ;
        RECT 721.010 795.720 724.770 796.690 ;
        RECT 725.610 795.720 728.450 796.690 ;
        RECT 729.290 795.720 733.050 796.690 ;
        RECT 733.890 795.720 737.650 796.690 ;
        RECT 738.490 795.720 741.330 796.690 ;
        RECT 742.170 795.720 745.930 796.690 ;
        RECT 746.770 795.720 750.530 796.690 ;
        RECT 751.370 795.720 754.210 796.690 ;
        RECT 755.050 795.720 758.810 796.690 ;
        RECT 759.650 795.720 763.410 796.690 ;
        RECT 764.250 795.720 767.090 796.690 ;
        RECT 767.930 795.720 771.690 796.690 ;
        RECT 772.530 795.720 776.290 796.690 ;
        RECT 777.130 795.720 779.970 796.690 ;
        RECT 780.810 795.720 784.570 796.690 ;
        RECT 785.410 795.720 789.170 796.690 ;
        RECT 790.010 795.720 792.850 796.690 ;
        RECT 793.690 795.720 797.450 796.690 ;
        RECT 0.100 4.280 798.000 795.720 ;
        RECT 0.650 0.155 3.490 4.280 ;
        RECT 4.330 0.155 8.090 4.280 ;
        RECT 8.930 0.155 12.690 4.280 ;
        RECT 13.530 0.155 16.370 4.280 ;
        RECT 17.210 0.155 20.970 4.280 ;
        RECT 21.810 0.155 25.570 4.280 ;
        RECT 26.410 0.155 29.250 4.280 ;
        RECT 30.090 0.155 33.850 4.280 ;
        RECT 34.690 0.155 38.450 4.280 ;
        RECT 39.290 0.155 42.130 4.280 ;
        RECT 42.970 0.155 46.730 4.280 ;
        RECT 47.570 0.155 51.330 4.280 ;
        RECT 52.170 0.155 55.010 4.280 ;
        RECT 55.850 0.155 59.610 4.280 ;
        RECT 60.450 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.890 4.280 ;
        RECT 68.730 0.155 72.490 4.280 ;
        RECT 73.330 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.770 4.280 ;
        RECT 81.610 0.155 85.370 4.280 ;
        RECT 86.210 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.650 4.280 ;
        RECT 94.490 0.155 98.250 4.280 ;
        RECT 99.090 0.155 102.850 4.280 ;
        RECT 103.690 0.155 107.450 4.280 ;
        RECT 108.290 0.155 111.130 4.280 ;
        RECT 111.970 0.155 115.730 4.280 ;
        RECT 116.570 0.155 120.330 4.280 ;
        RECT 121.170 0.155 124.010 4.280 ;
        RECT 124.850 0.155 128.610 4.280 ;
        RECT 129.450 0.155 133.210 4.280 ;
        RECT 134.050 0.155 136.890 4.280 ;
        RECT 137.730 0.155 141.490 4.280 ;
        RECT 142.330 0.155 146.090 4.280 ;
        RECT 146.930 0.155 149.770 4.280 ;
        RECT 150.610 0.155 154.370 4.280 ;
        RECT 155.210 0.155 158.970 4.280 ;
        RECT 159.810 0.155 162.650 4.280 ;
        RECT 163.490 0.155 167.250 4.280 ;
        RECT 168.090 0.155 171.850 4.280 ;
        RECT 172.690 0.155 175.530 4.280 ;
        RECT 176.370 0.155 180.130 4.280 ;
        RECT 180.970 0.155 184.730 4.280 ;
        RECT 185.570 0.155 188.410 4.280 ;
        RECT 189.250 0.155 193.010 4.280 ;
        RECT 193.850 0.155 197.610 4.280 ;
        RECT 198.450 0.155 201.290 4.280 ;
        RECT 202.130 0.155 205.890 4.280 ;
        RECT 206.730 0.155 210.490 4.280 ;
        RECT 211.330 0.155 215.090 4.280 ;
        RECT 215.930 0.155 218.770 4.280 ;
        RECT 219.610 0.155 223.370 4.280 ;
        RECT 224.210 0.155 227.970 4.280 ;
        RECT 228.810 0.155 231.650 4.280 ;
        RECT 232.490 0.155 236.250 4.280 ;
        RECT 237.090 0.155 240.850 4.280 ;
        RECT 241.690 0.155 244.530 4.280 ;
        RECT 245.370 0.155 249.130 4.280 ;
        RECT 249.970 0.155 253.730 4.280 ;
        RECT 254.570 0.155 257.410 4.280 ;
        RECT 258.250 0.155 262.010 4.280 ;
        RECT 262.850 0.155 266.610 4.280 ;
        RECT 267.450 0.155 270.290 4.280 ;
        RECT 271.130 0.155 274.890 4.280 ;
        RECT 275.730 0.155 279.490 4.280 ;
        RECT 280.330 0.155 283.170 4.280 ;
        RECT 284.010 0.155 287.770 4.280 ;
        RECT 288.610 0.155 292.370 4.280 ;
        RECT 293.210 0.155 296.050 4.280 ;
        RECT 296.890 0.155 300.650 4.280 ;
        RECT 301.490 0.155 305.250 4.280 ;
        RECT 306.090 0.155 309.850 4.280 ;
        RECT 310.690 0.155 313.530 4.280 ;
        RECT 314.370 0.155 318.130 4.280 ;
        RECT 318.970 0.155 322.730 4.280 ;
        RECT 323.570 0.155 326.410 4.280 ;
        RECT 327.250 0.155 331.010 4.280 ;
        RECT 331.850 0.155 335.610 4.280 ;
        RECT 336.450 0.155 339.290 4.280 ;
        RECT 340.130 0.155 343.890 4.280 ;
        RECT 344.730 0.155 348.490 4.280 ;
        RECT 349.330 0.155 352.170 4.280 ;
        RECT 353.010 0.155 356.770 4.280 ;
        RECT 357.610 0.155 361.370 4.280 ;
        RECT 362.210 0.155 365.050 4.280 ;
        RECT 365.890 0.155 369.650 4.280 ;
        RECT 370.490 0.155 374.250 4.280 ;
        RECT 375.090 0.155 377.930 4.280 ;
        RECT 378.770 0.155 382.530 4.280 ;
        RECT 383.370 0.155 387.130 4.280 ;
        RECT 387.970 0.155 390.810 4.280 ;
        RECT 391.650 0.155 395.410 4.280 ;
        RECT 396.250 0.155 400.010 4.280 ;
        RECT 400.850 0.155 403.690 4.280 ;
        RECT 404.530 0.155 408.290 4.280 ;
        RECT 409.130 0.155 412.890 4.280 ;
        RECT 413.730 0.155 417.490 4.280 ;
        RECT 418.330 0.155 421.170 4.280 ;
        RECT 422.010 0.155 425.770 4.280 ;
        RECT 426.610 0.155 430.370 4.280 ;
        RECT 431.210 0.155 434.050 4.280 ;
        RECT 434.890 0.155 438.650 4.280 ;
        RECT 439.490 0.155 443.250 4.280 ;
        RECT 444.090 0.155 446.930 4.280 ;
        RECT 447.770 0.155 451.530 4.280 ;
        RECT 452.370 0.155 456.130 4.280 ;
        RECT 456.970 0.155 459.810 4.280 ;
        RECT 460.650 0.155 464.410 4.280 ;
        RECT 465.250 0.155 469.010 4.280 ;
        RECT 469.850 0.155 472.690 4.280 ;
        RECT 473.530 0.155 477.290 4.280 ;
        RECT 478.130 0.155 481.890 4.280 ;
        RECT 482.730 0.155 485.570 4.280 ;
        RECT 486.410 0.155 490.170 4.280 ;
        RECT 491.010 0.155 494.770 4.280 ;
        RECT 495.610 0.155 498.450 4.280 ;
        RECT 499.290 0.155 503.050 4.280 ;
        RECT 503.890 0.155 507.650 4.280 ;
        RECT 508.490 0.155 511.330 4.280 ;
        RECT 512.170 0.155 515.930 4.280 ;
        RECT 516.770 0.155 520.530 4.280 ;
        RECT 521.370 0.155 525.130 4.280 ;
        RECT 525.970 0.155 528.810 4.280 ;
        RECT 529.650 0.155 533.410 4.280 ;
        RECT 534.250 0.155 538.010 4.280 ;
        RECT 538.850 0.155 541.690 4.280 ;
        RECT 542.530 0.155 546.290 4.280 ;
        RECT 547.130 0.155 550.890 4.280 ;
        RECT 551.730 0.155 554.570 4.280 ;
        RECT 555.410 0.155 559.170 4.280 ;
        RECT 560.010 0.155 563.770 4.280 ;
        RECT 564.610 0.155 567.450 4.280 ;
        RECT 568.290 0.155 572.050 4.280 ;
        RECT 572.890 0.155 576.650 4.280 ;
        RECT 577.490 0.155 580.330 4.280 ;
        RECT 581.170 0.155 584.930 4.280 ;
        RECT 585.770 0.155 589.530 4.280 ;
        RECT 590.370 0.155 593.210 4.280 ;
        RECT 594.050 0.155 597.810 4.280 ;
        RECT 598.650 0.155 602.410 4.280 ;
        RECT 603.250 0.155 606.090 4.280 ;
        RECT 606.930 0.155 610.690 4.280 ;
        RECT 611.530 0.155 615.290 4.280 ;
        RECT 616.130 0.155 619.890 4.280 ;
        RECT 620.730 0.155 623.570 4.280 ;
        RECT 624.410 0.155 628.170 4.280 ;
        RECT 629.010 0.155 632.770 4.280 ;
        RECT 633.610 0.155 636.450 4.280 ;
        RECT 637.290 0.155 641.050 4.280 ;
        RECT 641.890 0.155 645.650 4.280 ;
        RECT 646.490 0.155 649.330 4.280 ;
        RECT 650.170 0.155 653.930 4.280 ;
        RECT 654.770 0.155 658.530 4.280 ;
        RECT 659.370 0.155 662.210 4.280 ;
        RECT 663.050 0.155 666.810 4.280 ;
        RECT 667.650 0.155 671.410 4.280 ;
        RECT 672.250 0.155 675.090 4.280 ;
        RECT 675.930 0.155 679.690 4.280 ;
        RECT 680.530 0.155 684.290 4.280 ;
        RECT 685.130 0.155 687.970 4.280 ;
        RECT 688.810 0.155 692.570 4.280 ;
        RECT 693.410 0.155 697.170 4.280 ;
        RECT 698.010 0.155 700.850 4.280 ;
        RECT 701.690 0.155 705.450 4.280 ;
        RECT 706.290 0.155 710.050 4.280 ;
        RECT 710.890 0.155 713.730 4.280 ;
        RECT 714.570 0.155 718.330 4.280 ;
        RECT 719.170 0.155 722.930 4.280 ;
        RECT 723.770 0.155 727.530 4.280 ;
        RECT 728.370 0.155 731.210 4.280 ;
        RECT 732.050 0.155 735.810 4.280 ;
        RECT 736.650 0.155 740.410 4.280 ;
        RECT 741.250 0.155 744.090 4.280 ;
        RECT 744.930 0.155 748.690 4.280 ;
        RECT 749.530 0.155 753.290 4.280 ;
        RECT 754.130 0.155 756.970 4.280 ;
        RECT 757.810 0.155 761.570 4.280 ;
        RECT 762.410 0.155 766.170 4.280 ;
        RECT 767.010 0.155 769.850 4.280 ;
        RECT 770.690 0.155 774.450 4.280 ;
        RECT 775.290 0.155 779.050 4.280 ;
        RECT 779.890 0.155 782.730 4.280 ;
        RECT 783.570 0.155 787.330 4.280 ;
        RECT 788.170 0.155 791.930 4.280 ;
        RECT 792.770 0.155 795.610 4.280 ;
        RECT 796.450 0.155 798.000 4.280 ;
      LAYER met3 ;
        RECT 4.400 795.240 795.600 796.105 ;
        RECT 4.000 789.840 796.000 795.240 ;
        RECT 4.400 788.440 795.600 789.840 ;
        RECT 4.000 784.400 796.000 788.440 ;
        RECT 4.000 783.040 795.600 784.400 ;
        RECT 4.400 783.000 795.600 783.040 ;
        RECT 4.400 781.640 796.000 783.000 ;
        RECT 4.000 777.600 796.000 781.640 ;
        RECT 4.400 776.200 795.600 777.600 ;
        RECT 4.000 770.800 796.000 776.200 ;
        RECT 4.400 769.400 795.600 770.800 ;
        RECT 4.000 765.360 796.000 769.400 ;
        RECT 4.000 764.000 795.600 765.360 ;
        RECT 4.400 763.960 795.600 764.000 ;
        RECT 4.400 762.600 796.000 763.960 ;
        RECT 4.000 758.560 796.000 762.600 ;
        RECT 4.000 757.200 795.600 758.560 ;
        RECT 4.400 757.160 795.600 757.200 ;
        RECT 4.400 755.800 796.000 757.160 ;
        RECT 4.000 751.760 796.000 755.800 ;
        RECT 4.400 750.360 795.600 751.760 ;
        RECT 4.000 746.320 796.000 750.360 ;
        RECT 4.000 744.960 795.600 746.320 ;
        RECT 4.400 744.920 795.600 744.960 ;
        RECT 4.400 743.560 796.000 744.920 ;
        RECT 4.000 739.520 796.000 743.560 ;
        RECT 4.000 738.160 795.600 739.520 ;
        RECT 4.400 738.120 795.600 738.160 ;
        RECT 4.400 736.760 796.000 738.120 ;
        RECT 4.000 732.720 796.000 736.760 ;
        RECT 4.400 731.320 795.600 732.720 ;
        RECT 4.000 727.280 796.000 731.320 ;
        RECT 4.000 725.920 795.600 727.280 ;
        RECT 4.400 725.880 795.600 725.920 ;
        RECT 4.400 724.520 796.000 725.880 ;
        RECT 4.000 720.480 796.000 724.520 ;
        RECT 4.000 719.120 795.600 720.480 ;
        RECT 4.400 719.080 795.600 719.120 ;
        RECT 4.400 717.720 796.000 719.080 ;
        RECT 4.000 713.680 796.000 717.720 ;
        RECT 4.400 712.280 795.600 713.680 ;
        RECT 4.000 708.240 796.000 712.280 ;
        RECT 4.000 706.880 795.600 708.240 ;
        RECT 4.400 706.840 795.600 706.880 ;
        RECT 4.400 705.480 796.000 706.840 ;
        RECT 4.000 701.440 796.000 705.480 ;
        RECT 4.000 700.080 795.600 701.440 ;
        RECT 4.400 700.040 795.600 700.080 ;
        RECT 4.400 698.680 796.000 700.040 ;
        RECT 4.000 694.640 796.000 698.680 ;
        RECT 4.400 693.240 795.600 694.640 ;
        RECT 4.000 689.200 796.000 693.240 ;
        RECT 4.000 687.840 795.600 689.200 ;
        RECT 4.400 687.800 795.600 687.840 ;
        RECT 4.400 686.440 796.000 687.800 ;
        RECT 4.000 682.400 796.000 686.440 ;
        RECT 4.000 681.040 795.600 682.400 ;
        RECT 4.400 681.000 795.600 681.040 ;
        RECT 4.400 679.640 796.000 681.000 ;
        RECT 4.000 675.600 796.000 679.640 ;
        RECT 4.400 674.200 795.600 675.600 ;
        RECT 4.000 670.160 796.000 674.200 ;
        RECT 4.000 668.800 795.600 670.160 ;
        RECT 4.400 668.760 795.600 668.800 ;
        RECT 4.400 667.400 796.000 668.760 ;
        RECT 4.000 663.360 796.000 667.400 ;
        RECT 4.000 662.000 795.600 663.360 ;
        RECT 4.400 661.960 795.600 662.000 ;
        RECT 4.400 660.600 796.000 661.960 ;
        RECT 4.000 656.560 796.000 660.600 ;
        RECT 4.400 655.160 795.600 656.560 ;
        RECT 4.000 651.120 796.000 655.160 ;
        RECT 4.000 649.760 795.600 651.120 ;
        RECT 4.400 649.720 795.600 649.760 ;
        RECT 4.400 648.360 796.000 649.720 ;
        RECT 4.000 644.320 796.000 648.360 ;
        RECT 4.000 642.960 795.600 644.320 ;
        RECT 4.400 642.920 795.600 642.960 ;
        RECT 4.400 641.560 796.000 642.920 ;
        RECT 4.000 637.520 796.000 641.560 ;
        RECT 4.400 636.120 795.600 637.520 ;
        RECT 4.000 630.720 796.000 636.120 ;
        RECT 4.400 629.320 795.600 630.720 ;
        RECT 4.000 625.280 796.000 629.320 ;
        RECT 4.000 623.920 795.600 625.280 ;
        RECT 4.400 623.880 795.600 623.920 ;
        RECT 4.400 622.520 796.000 623.880 ;
        RECT 4.000 618.480 796.000 622.520 ;
        RECT 4.400 617.080 795.600 618.480 ;
        RECT 4.000 611.680 796.000 617.080 ;
        RECT 4.400 610.280 795.600 611.680 ;
        RECT 4.000 606.240 796.000 610.280 ;
        RECT 4.000 604.880 795.600 606.240 ;
        RECT 4.400 604.840 795.600 604.880 ;
        RECT 4.400 603.480 796.000 604.840 ;
        RECT 4.000 599.440 796.000 603.480 ;
        RECT 4.000 598.080 795.600 599.440 ;
        RECT 4.400 598.040 795.600 598.080 ;
        RECT 4.400 596.680 796.000 598.040 ;
        RECT 4.000 592.640 796.000 596.680 ;
        RECT 4.400 591.240 795.600 592.640 ;
        RECT 4.000 587.200 796.000 591.240 ;
        RECT 4.000 585.840 795.600 587.200 ;
        RECT 4.400 585.800 795.600 585.840 ;
        RECT 4.400 584.440 796.000 585.800 ;
        RECT 4.000 580.400 796.000 584.440 ;
        RECT 4.000 579.040 795.600 580.400 ;
        RECT 4.400 579.000 795.600 579.040 ;
        RECT 4.400 577.640 796.000 579.000 ;
        RECT 4.000 573.600 796.000 577.640 ;
        RECT 4.400 572.200 795.600 573.600 ;
        RECT 4.000 568.160 796.000 572.200 ;
        RECT 4.000 566.800 795.600 568.160 ;
        RECT 4.400 566.760 795.600 566.800 ;
        RECT 4.400 565.400 796.000 566.760 ;
        RECT 4.000 561.360 796.000 565.400 ;
        RECT 4.000 560.000 795.600 561.360 ;
        RECT 4.400 559.960 795.600 560.000 ;
        RECT 4.400 558.600 796.000 559.960 ;
        RECT 4.000 554.560 796.000 558.600 ;
        RECT 4.400 553.160 795.600 554.560 ;
        RECT 4.000 549.120 796.000 553.160 ;
        RECT 4.000 547.760 795.600 549.120 ;
        RECT 4.400 547.720 795.600 547.760 ;
        RECT 4.400 546.360 796.000 547.720 ;
        RECT 4.000 542.320 796.000 546.360 ;
        RECT 4.000 540.960 795.600 542.320 ;
        RECT 4.400 540.920 795.600 540.960 ;
        RECT 4.400 539.560 796.000 540.920 ;
        RECT 4.000 535.520 796.000 539.560 ;
        RECT 4.400 534.120 795.600 535.520 ;
        RECT 4.000 530.080 796.000 534.120 ;
        RECT 4.000 528.720 795.600 530.080 ;
        RECT 4.400 528.680 795.600 528.720 ;
        RECT 4.400 527.320 796.000 528.680 ;
        RECT 4.000 523.280 796.000 527.320 ;
        RECT 4.000 521.920 795.600 523.280 ;
        RECT 4.400 521.880 795.600 521.920 ;
        RECT 4.400 520.520 796.000 521.880 ;
        RECT 4.000 516.480 796.000 520.520 ;
        RECT 4.400 515.080 795.600 516.480 ;
        RECT 4.000 511.040 796.000 515.080 ;
        RECT 4.000 509.680 795.600 511.040 ;
        RECT 4.400 509.640 795.600 509.680 ;
        RECT 4.400 508.280 796.000 509.640 ;
        RECT 4.000 504.240 796.000 508.280 ;
        RECT 4.000 502.880 795.600 504.240 ;
        RECT 4.400 502.840 795.600 502.880 ;
        RECT 4.400 501.480 796.000 502.840 ;
        RECT 4.000 497.440 796.000 501.480 ;
        RECT 4.400 496.040 795.600 497.440 ;
        RECT 4.000 490.640 796.000 496.040 ;
        RECT 4.400 489.240 795.600 490.640 ;
        RECT 4.000 485.200 796.000 489.240 ;
        RECT 4.000 483.840 795.600 485.200 ;
        RECT 4.400 483.800 795.600 483.840 ;
        RECT 4.400 482.440 796.000 483.800 ;
        RECT 4.000 478.400 796.000 482.440 ;
        RECT 4.400 477.000 795.600 478.400 ;
        RECT 4.000 471.600 796.000 477.000 ;
        RECT 4.400 470.200 795.600 471.600 ;
        RECT 4.000 466.160 796.000 470.200 ;
        RECT 4.000 464.800 795.600 466.160 ;
        RECT 4.400 464.760 795.600 464.800 ;
        RECT 4.400 463.400 796.000 464.760 ;
        RECT 4.000 459.360 796.000 463.400 ;
        RECT 4.400 457.960 795.600 459.360 ;
        RECT 4.000 452.560 796.000 457.960 ;
        RECT 4.400 451.160 795.600 452.560 ;
        RECT 4.000 447.120 796.000 451.160 ;
        RECT 4.000 445.760 795.600 447.120 ;
        RECT 4.400 445.720 795.600 445.760 ;
        RECT 4.400 444.360 796.000 445.720 ;
        RECT 4.000 440.320 796.000 444.360 ;
        RECT 4.000 438.960 795.600 440.320 ;
        RECT 4.400 438.920 795.600 438.960 ;
        RECT 4.400 437.560 796.000 438.920 ;
        RECT 4.000 433.520 796.000 437.560 ;
        RECT 4.400 432.120 795.600 433.520 ;
        RECT 4.000 428.080 796.000 432.120 ;
        RECT 4.000 426.720 795.600 428.080 ;
        RECT 4.400 426.680 795.600 426.720 ;
        RECT 4.400 425.320 796.000 426.680 ;
        RECT 4.000 421.280 796.000 425.320 ;
        RECT 4.000 419.920 795.600 421.280 ;
        RECT 4.400 419.880 795.600 419.920 ;
        RECT 4.400 418.520 796.000 419.880 ;
        RECT 4.000 414.480 796.000 418.520 ;
        RECT 4.400 413.080 795.600 414.480 ;
        RECT 4.000 409.040 796.000 413.080 ;
        RECT 4.000 407.680 795.600 409.040 ;
        RECT 4.400 407.640 795.600 407.680 ;
        RECT 4.400 406.280 796.000 407.640 ;
        RECT 4.000 402.240 796.000 406.280 ;
        RECT 4.000 400.880 795.600 402.240 ;
        RECT 4.400 400.840 795.600 400.880 ;
        RECT 4.400 399.480 796.000 400.840 ;
        RECT 4.000 395.440 796.000 399.480 ;
        RECT 4.400 394.040 795.600 395.440 ;
        RECT 4.000 390.000 796.000 394.040 ;
        RECT 4.000 388.640 795.600 390.000 ;
        RECT 4.400 388.600 795.600 388.640 ;
        RECT 4.400 387.240 796.000 388.600 ;
        RECT 4.000 383.200 796.000 387.240 ;
        RECT 4.000 381.840 795.600 383.200 ;
        RECT 4.400 381.800 795.600 381.840 ;
        RECT 4.400 380.440 796.000 381.800 ;
        RECT 4.000 376.400 796.000 380.440 ;
        RECT 4.400 375.000 795.600 376.400 ;
        RECT 4.000 370.960 796.000 375.000 ;
        RECT 4.000 369.600 795.600 370.960 ;
        RECT 4.400 369.560 795.600 369.600 ;
        RECT 4.400 368.200 796.000 369.560 ;
        RECT 4.000 364.160 796.000 368.200 ;
        RECT 4.000 362.800 795.600 364.160 ;
        RECT 4.400 362.760 795.600 362.800 ;
        RECT 4.400 361.400 796.000 362.760 ;
        RECT 4.000 357.360 796.000 361.400 ;
        RECT 4.400 355.960 795.600 357.360 ;
        RECT 4.000 351.920 796.000 355.960 ;
        RECT 4.000 350.560 795.600 351.920 ;
        RECT 4.400 350.520 795.600 350.560 ;
        RECT 4.400 349.160 796.000 350.520 ;
        RECT 4.000 345.120 796.000 349.160 ;
        RECT 4.000 343.760 795.600 345.120 ;
        RECT 4.400 343.720 795.600 343.760 ;
        RECT 4.400 342.360 796.000 343.720 ;
        RECT 4.000 338.320 796.000 342.360 ;
        RECT 4.400 336.920 795.600 338.320 ;
        RECT 4.000 331.520 796.000 336.920 ;
        RECT 4.400 330.120 795.600 331.520 ;
        RECT 4.000 326.080 796.000 330.120 ;
        RECT 4.000 324.720 795.600 326.080 ;
        RECT 4.400 324.680 795.600 324.720 ;
        RECT 4.400 323.320 796.000 324.680 ;
        RECT 4.000 319.280 796.000 323.320 ;
        RECT 4.400 317.880 795.600 319.280 ;
        RECT 4.000 312.480 796.000 317.880 ;
        RECT 4.400 311.080 795.600 312.480 ;
        RECT 4.000 307.040 796.000 311.080 ;
        RECT 4.000 305.680 795.600 307.040 ;
        RECT 4.400 305.640 795.600 305.680 ;
        RECT 4.400 304.280 796.000 305.640 ;
        RECT 4.000 300.240 796.000 304.280 ;
        RECT 4.000 298.880 795.600 300.240 ;
        RECT 4.400 298.840 795.600 298.880 ;
        RECT 4.400 297.480 796.000 298.840 ;
        RECT 4.000 293.440 796.000 297.480 ;
        RECT 4.400 292.040 795.600 293.440 ;
        RECT 4.000 288.000 796.000 292.040 ;
        RECT 4.000 286.640 795.600 288.000 ;
        RECT 4.400 286.600 795.600 286.640 ;
        RECT 4.400 285.240 796.000 286.600 ;
        RECT 4.000 281.200 796.000 285.240 ;
        RECT 4.000 279.840 795.600 281.200 ;
        RECT 4.400 279.800 795.600 279.840 ;
        RECT 4.400 278.440 796.000 279.800 ;
        RECT 4.000 274.400 796.000 278.440 ;
        RECT 4.400 273.000 795.600 274.400 ;
        RECT 4.000 268.960 796.000 273.000 ;
        RECT 4.000 267.600 795.600 268.960 ;
        RECT 4.400 267.560 795.600 267.600 ;
        RECT 4.400 266.200 796.000 267.560 ;
        RECT 4.000 262.160 796.000 266.200 ;
        RECT 4.000 260.800 795.600 262.160 ;
        RECT 4.400 260.760 795.600 260.800 ;
        RECT 4.400 259.400 796.000 260.760 ;
        RECT 4.000 255.360 796.000 259.400 ;
        RECT 4.400 253.960 795.600 255.360 ;
        RECT 4.000 249.920 796.000 253.960 ;
        RECT 4.000 248.560 795.600 249.920 ;
        RECT 4.400 248.520 795.600 248.560 ;
        RECT 4.400 247.160 796.000 248.520 ;
        RECT 4.000 243.120 796.000 247.160 ;
        RECT 4.000 241.760 795.600 243.120 ;
        RECT 4.400 241.720 795.600 241.760 ;
        RECT 4.400 240.360 796.000 241.720 ;
        RECT 4.000 236.320 796.000 240.360 ;
        RECT 4.400 234.920 795.600 236.320 ;
        RECT 4.000 230.880 796.000 234.920 ;
        RECT 4.000 229.520 795.600 230.880 ;
        RECT 4.400 229.480 795.600 229.520 ;
        RECT 4.400 228.120 796.000 229.480 ;
        RECT 4.000 224.080 796.000 228.120 ;
        RECT 4.000 222.720 795.600 224.080 ;
        RECT 4.400 222.680 795.600 222.720 ;
        RECT 4.400 221.320 796.000 222.680 ;
        RECT 4.000 217.280 796.000 221.320 ;
        RECT 4.400 215.880 795.600 217.280 ;
        RECT 4.000 211.840 796.000 215.880 ;
        RECT 4.000 210.480 795.600 211.840 ;
        RECT 4.400 210.440 795.600 210.480 ;
        RECT 4.400 209.080 796.000 210.440 ;
        RECT 4.000 205.040 796.000 209.080 ;
        RECT 4.000 203.680 795.600 205.040 ;
        RECT 4.400 203.640 795.600 203.680 ;
        RECT 4.400 202.280 796.000 203.640 ;
        RECT 4.000 198.240 796.000 202.280 ;
        RECT 4.400 196.840 795.600 198.240 ;
        RECT 4.000 192.800 796.000 196.840 ;
        RECT 4.000 191.440 795.600 192.800 ;
        RECT 4.400 191.400 795.600 191.440 ;
        RECT 4.400 190.040 796.000 191.400 ;
        RECT 4.000 186.000 796.000 190.040 ;
        RECT 4.000 184.640 795.600 186.000 ;
        RECT 4.400 184.600 795.600 184.640 ;
        RECT 4.400 183.240 796.000 184.600 ;
        RECT 4.000 179.200 796.000 183.240 ;
        RECT 4.400 177.800 795.600 179.200 ;
        RECT 4.000 172.400 796.000 177.800 ;
        RECT 4.400 171.000 795.600 172.400 ;
        RECT 4.000 166.960 796.000 171.000 ;
        RECT 4.000 165.600 795.600 166.960 ;
        RECT 4.400 165.560 795.600 165.600 ;
        RECT 4.400 164.200 796.000 165.560 ;
        RECT 4.000 160.160 796.000 164.200 ;
        RECT 4.400 158.760 795.600 160.160 ;
        RECT 4.000 153.360 796.000 158.760 ;
        RECT 4.400 151.960 795.600 153.360 ;
        RECT 4.000 147.920 796.000 151.960 ;
        RECT 4.000 146.560 795.600 147.920 ;
        RECT 4.400 146.520 795.600 146.560 ;
        RECT 4.400 145.160 796.000 146.520 ;
        RECT 4.000 141.120 796.000 145.160 ;
        RECT 4.000 139.760 795.600 141.120 ;
        RECT 4.400 139.720 795.600 139.760 ;
        RECT 4.400 138.360 796.000 139.720 ;
        RECT 4.000 134.320 796.000 138.360 ;
        RECT 4.400 132.920 795.600 134.320 ;
        RECT 4.000 128.880 796.000 132.920 ;
        RECT 4.000 127.520 795.600 128.880 ;
        RECT 4.400 127.480 795.600 127.520 ;
        RECT 4.400 126.120 796.000 127.480 ;
        RECT 4.000 122.080 796.000 126.120 ;
        RECT 4.000 120.720 795.600 122.080 ;
        RECT 4.400 120.680 795.600 120.720 ;
        RECT 4.400 119.320 796.000 120.680 ;
        RECT 4.000 115.280 796.000 119.320 ;
        RECT 4.400 113.880 795.600 115.280 ;
        RECT 4.000 109.840 796.000 113.880 ;
        RECT 4.000 108.480 795.600 109.840 ;
        RECT 4.400 108.440 795.600 108.480 ;
        RECT 4.400 107.080 796.000 108.440 ;
        RECT 4.000 103.040 796.000 107.080 ;
        RECT 4.000 101.680 795.600 103.040 ;
        RECT 4.400 101.640 795.600 101.680 ;
        RECT 4.400 100.280 796.000 101.640 ;
        RECT 4.000 96.240 796.000 100.280 ;
        RECT 4.400 94.840 795.600 96.240 ;
        RECT 4.000 90.800 796.000 94.840 ;
        RECT 4.000 89.440 795.600 90.800 ;
        RECT 4.400 89.400 795.600 89.440 ;
        RECT 4.400 88.040 796.000 89.400 ;
        RECT 4.000 84.000 796.000 88.040 ;
        RECT 4.000 82.640 795.600 84.000 ;
        RECT 4.400 82.600 795.600 82.640 ;
        RECT 4.400 81.240 796.000 82.600 ;
        RECT 4.000 77.200 796.000 81.240 ;
        RECT 4.400 75.800 795.600 77.200 ;
        RECT 4.000 71.760 796.000 75.800 ;
        RECT 4.000 70.400 795.600 71.760 ;
        RECT 4.400 70.360 795.600 70.400 ;
        RECT 4.400 69.000 796.000 70.360 ;
        RECT 4.000 64.960 796.000 69.000 ;
        RECT 4.000 63.600 795.600 64.960 ;
        RECT 4.400 63.560 795.600 63.600 ;
        RECT 4.400 62.200 796.000 63.560 ;
        RECT 4.000 58.160 796.000 62.200 ;
        RECT 4.400 56.760 795.600 58.160 ;
        RECT 4.000 52.720 796.000 56.760 ;
        RECT 4.000 51.360 795.600 52.720 ;
        RECT 4.400 51.320 795.600 51.360 ;
        RECT 4.400 49.960 796.000 51.320 ;
        RECT 4.000 45.920 796.000 49.960 ;
        RECT 4.000 44.560 795.600 45.920 ;
        RECT 4.400 44.520 795.600 44.560 ;
        RECT 4.400 43.160 796.000 44.520 ;
        RECT 4.000 39.120 796.000 43.160 ;
        RECT 4.400 37.720 795.600 39.120 ;
        RECT 4.000 32.320 796.000 37.720 ;
        RECT 4.400 30.920 795.600 32.320 ;
        RECT 4.000 26.880 796.000 30.920 ;
        RECT 4.000 25.520 795.600 26.880 ;
        RECT 4.400 25.480 795.600 25.520 ;
        RECT 4.400 24.120 796.000 25.480 ;
        RECT 4.000 20.080 796.000 24.120 ;
        RECT 4.400 18.680 795.600 20.080 ;
        RECT 4.000 13.280 796.000 18.680 ;
        RECT 4.400 11.880 795.600 13.280 ;
        RECT 4.000 7.840 796.000 11.880 ;
        RECT 4.000 6.480 795.600 7.840 ;
        RECT 4.400 6.440 795.600 6.480 ;
        RECT 4.400 5.080 796.000 6.440 ;
        RECT 4.000 1.040 796.000 5.080 ;
        RECT 4.000 0.175 795.600 1.040 ;
      LAYER met4 ;
        RECT 352.655 38.935 404.640 621.345 ;
        RECT 407.040 38.935 481.440 621.345 ;
        RECT 483.840 38.935 558.240 621.345 ;
        RECT 560.640 38.935 635.040 621.345 ;
        RECT 637.440 38.935 711.840 621.345 ;
        RECT 714.240 38.935 785.385 621.345 ;
  END
END MEM_WB
END LIBRARY

