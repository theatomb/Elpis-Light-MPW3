VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO custom_sram
  CLASS BLOCK ;
  FOREIGN custom_sram ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 1500.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 26.560 1800.000 27.160 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 1496.000 637.470 1500.000 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 1496.000 937.390 1500.000 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 0.000 956.250 4.000 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 615.440 1800.000 616.040 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 722.880 1800.000 723.480 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.960 4.000 1237.560 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 937.080 1800.000 937.680 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 133.320 1800.000 133.920 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 240.760 1800.000 241.360 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 293.800 1800.000 294.400 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 1496.000 187.590 1500.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.200 4.000 637.800 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 1496.000 337.550 1500.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 454.960 1800.000 455.560 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 1496.000 412.530 1500.000 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 1496.000 487.510 1500.000 ;
    END
  END a[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END clk
  PIN csb0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END csb0_to_sram
  PIN d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 1496.000 37.630 1500.000 ;
    END
  END d[0]
  PIN d[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END d[10]
  PIN d[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 1496.000 712.450 1500.000 ;
    END
  END d[11]
  PIN d[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 1496.000 787.430 1500.000 ;
    END
  END d[12]
  PIN d[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1087.360 4.000 1087.960 ;
    END
  END d[13]
  PIN d[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.160 4.000 1162.760 ;
    END
  END d[14]
  PIN d[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.670 0.000 1068.950 4.000 ;
    END
  END d[15]
  PIN d[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 669.160 1800.000 669.760 ;
    END
  END d[16]
  PIN d[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 776.600 1800.000 777.200 ;
    END
  END d[17]
  PIN d[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 883.360 1800.000 883.960 ;
    END
  END d[18]
  PIN d[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.610 0.000 1293.890 4.000 ;
    END
  END d[19]
  PIN d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 1496.000 112.610 1500.000 ;
    END
  END d[1]
  PIN d[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1312.440 4.000 1313.040 ;
    END
  END d[20]
  PIN d[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.010 1496.000 1312.290 1500.000 ;
    END
  END d[21]
  PIN d[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 1496.000 1462.250 1500.000 ;
    END
  END d[22]
  PIN d[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1097.560 1800.000 1098.160 ;
    END
  END d[23]
  PIN d[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.950 1496.000 1537.230 1500.000 ;
    END
  END d[24]
  PIN d[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.930 1496.000 1612.210 1500.000 ;
    END
  END d[25]
  PIN d[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1205.000 1800.000 1205.600 ;
    END
  END d[26]
  PIN d[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.910 1496.000 1687.190 1500.000 ;
    END
  END d[27]
  PIN d[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.890 1496.000 1762.170 1500.000 ;
    END
  END d[28]
  PIN d[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1311.760 1800.000 1312.360 ;
    END
  END d[29]
  PIN d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END d[2]
  PIN d[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.790 0.000 1631.070 4.000 ;
    END
  END d[30]
  PIN d[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1472.920 1800.000 1473.520 ;
    END
  END d[31]
  PIN d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 347.520 1800.000 348.120 ;
    END
  END d[3]
  PIN d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 401.240 1800.000 401.840 ;
    END
  END d[4]
  PIN d[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 1496.000 262.570 1500.000 ;
    END
  END d[5]
  PIN d[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.000 4.000 712.600 ;
    END
  END d[6]
  PIN d[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END d[7]
  PIN d[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END d[8]
  PIN d[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 508.680 1800.000 509.280 ;
    END
  END d[9]
  PIN q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 79.600 1800.000 80.200 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.080 4.000 937.680 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END q[11]
  PIN q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 1496.000 862.410 1500.000 ;
    END
  END q[12]
  PIN q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 561.720 1800.000 562.320 ;
    END
  END q[13]
  PIN q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.090 1496.000 1012.370 1500.000 ;
    END
  END q[14]
  PIN q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.070 1496.000 1087.350 1500.000 ;
    END
  END q[15]
  PIN q[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 1496.000 1162.330 1500.000 ;
    END
  END q[16]
  PIN q[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 829.640 1800.000 830.240 ;
    END
  END q[17]
  PIN q[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END q[18]
  PIN q[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 990.800 1800.000 991.400 ;
    END
  END q[19]
  PIN q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 187.040 1800.000 187.640 ;
    END
  END q[1]
  PIN q[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030 1496.000 1237.310 1500.000 ;
    END
  END q[20]
  PIN q[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.990 1496.000 1387.270 1500.000 ;
    END
  END q[21]
  PIN q[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1043.840 1800.000 1044.440 ;
    END
  END q[22]
  PIN q[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 0.000 1406.130 4.000 ;
    END
  END q[23]
  PIN q[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.550 0.000 1518.830 4.000 ;
    END
  END q[24]
  PIN q[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1151.280 1800.000 1151.880 ;
    END
  END q[25]
  PIN q[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1387.240 4.000 1387.840 ;
    END
  END q[26]
  PIN q[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1258.720 1800.000 1259.320 ;
    END
  END q[27]
  PIN q[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END q[28]
  PIN q[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1365.480 1800.000 1366.080 ;
    END
  END q[29]
  PIN q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END q[2]
  PIN q[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1419.200 1800.000 1419.800 ;
    END
  END q[30]
  PIN q[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.490 0.000 1743.770 4.000 ;
    END
  END q[31]
  PIN q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 1496.000 562.490 1500.000 ;
    END
  END q[9]
  PIN spare_wen0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1488.080 ;
    END
  END vssd1
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END we
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1796.615 1487.925 ;
      LAYER met1 ;
        RECT 5.520 9.220 1796.675 1488.480 ;
      LAYER met2 ;
        RECT 6.990 1495.720 37.070 1496.410 ;
        RECT 37.910 1495.720 112.050 1496.410 ;
        RECT 112.890 1495.720 187.030 1496.410 ;
        RECT 187.870 1495.720 262.010 1496.410 ;
        RECT 262.850 1495.720 336.990 1496.410 ;
        RECT 337.830 1495.720 411.970 1496.410 ;
        RECT 412.810 1495.720 486.950 1496.410 ;
        RECT 487.790 1495.720 561.930 1496.410 ;
        RECT 562.770 1495.720 636.910 1496.410 ;
        RECT 637.750 1495.720 711.890 1496.410 ;
        RECT 712.730 1495.720 786.870 1496.410 ;
        RECT 787.710 1495.720 861.850 1496.410 ;
        RECT 862.690 1495.720 936.830 1496.410 ;
        RECT 937.670 1495.720 1011.810 1496.410 ;
        RECT 1012.650 1495.720 1086.790 1496.410 ;
        RECT 1087.630 1495.720 1161.770 1496.410 ;
        RECT 1162.610 1495.720 1236.750 1496.410 ;
        RECT 1237.590 1495.720 1311.730 1496.410 ;
        RECT 1312.570 1495.720 1386.710 1496.410 ;
        RECT 1387.550 1495.720 1461.690 1496.410 ;
        RECT 1462.530 1495.720 1536.670 1496.410 ;
        RECT 1537.510 1495.720 1611.650 1496.410 ;
        RECT 1612.490 1495.720 1686.630 1496.410 ;
        RECT 1687.470 1495.720 1761.610 1496.410 ;
        RECT 1762.450 1495.720 1795.740 1496.410 ;
        RECT 6.990 4.280 1795.740 1495.720 ;
        RECT 6.990 4.000 55.930 4.280 ;
        RECT 56.770 4.000 168.170 4.280 ;
        RECT 169.010 4.000 280.870 4.280 ;
        RECT 281.710 4.000 393.110 4.280 ;
        RECT 393.950 4.000 505.810 4.280 ;
        RECT 506.650 4.000 618.050 4.280 ;
        RECT 618.890 4.000 730.750 4.280 ;
        RECT 731.590 4.000 842.990 4.280 ;
        RECT 843.830 4.000 955.690 4.280 ;
        RECT 956.530 4.000 1068.390 4.280 ;
        RECT 1069.230 4.000 1180.630 4.280 ;
        RECT 1181.470 4.000 1293.330 4.280 ;
        RECT 1294.170 4.000 1405.570 4.280 ;
        RECT 1406.410 4.000 1518.270 4.280 ;
        RECT 1519.110 4.000 1630.510 4.280 ;
        RECT 1631.350 4.000 1743.210 4.280 ;
        RECT 1744.050 4.000 1795.740 4.280 ;
      LAYER met3 ;
        RECT 4.000 1473.920 1796.000 1488.005 ;
        RECT 4.000 1472.520 1795.600 1473.920 ;
        RECT 4.000 1463.040 1796.000 1472.520 ;
        RECT 4.400 1461.640 1796.000 1463.040 ;
        RECT 4.000 1420.200 1796.000 1461.640 ;
        RECT 4.000 1418.800 1795.600 1420.200 ;
        RECT 4.000 1388.240 1796.000 1418.800 ;
        RECT 4.400 1386.840 1796.000 1388.240 ;
        RECT 4.000 1366.480 1796.000 1386.840 ;
        RECT 4.000 1365.080 1795.600 1366.480 ;
        RECT 4.000 1313.440 1796.000 1365.080 ;
        RECT 4.400 1312.760 1796.000 1313.440 ;
        RECT 4.400 1312.040 1795.600 1312.760 ;
        RECT 4.000 1311.360 1795.600 1312.040 ;
        RECT 4.000 1259.720 1796.000 1311.360 ;
        RECT 4.000 1258.320 1795.600 1259.720 ;
        RECT 4.000 1237.960 1796.000 1258.320 ;
        RECT 4.400 1236.560 1796.000 1237.960 ;
        RECT 4.000 1206.000 1796.000 1236.560 ;
        RECT 4.000 1204.600 1795.600 1206.000 ;
        RECT 4.000 1163.160 1796.000 1204.600 ;
        RECT 4.400 1161.760 1796.000 1163.160 ;
        RECT 4.000 1152.280 1796.000 1161.760 ;
        RECT 4.000 1150.880 1795.600 1152.280 ;
        RECT 4.000 1098.560 1796.000 1150.880 ;
        RECT 4.000 1097.160 1795.600 1098.560 ;
        RECT 4.000 1088.360 1796.000 1097.160 ;
        RECT 4.400 1086.960 1796.000 1088.360 ;
        RECT 4.000 1044.840 1796.000 1086.960 ;
        RECT 4.000 1043.440 1795.600 1044.840 ;
        RECT 4.000 1012.880 1796.000 1043.440 ;
        RECT 4.400 1011.480 1796.000 1012.880 ;
        RECT 4.000 991.800 1796.000 1011.480 ;
        RECT 4.000 990.400 1795.600 991.800 ;
        RECT 4.000 938.080 1796.000 990.400 ;
        RECT 4.400 936.680 1795.600 938.080 ;
        RECT 4.000 884.360 1796.000 936.680 ;
        RECT 4.000 882.960 1795.600 884.360 ;
        RECT 4.000 863.280 1796.000 882.960 ;
        RECT 4.400 861.880 1796.000 863.280 ;
        RECT 4.000 830.640 1796.000 861.880 ;
        RECT 4.000 829.240 1795.600 830.640 ;
        RECT 4.000 788.480 1796.000 829.240 ;
        RECT 4.400 787.080 1796.000 788.480 ;
        RECT 4.000 777.600 1796.000 787.080 ;
        RECT 4.000 776.200 1795.600 777.600 ;
        RECT 4.000 723.880 1796.000 776.200 ;
        RECT 4.000 722.480 1795.600 723.880 ;
        RECT 4.000 713.000 1796.000 722.480 ;
        RECT 4.400 711.600 1796.000 713.000 ;
        RECT 4.000 670.160 1796.000 711.600 ;
        RECT 4.000 668.760 1795.600 670.160 ;
        RECT 4.000 638.200 1796.000 668.760 ;
        RECT 4.400 636.800 1796.000 638.200 ;
        RECT 4.000 616.440 1796.000 636.800 ;
        RECT 4.000 615.040 1795.600 616.440 ;
        RECT 4.000 563.400 1796.000 615.040 ;
        RECT 4.400 562.720 1796.000 563.400 ;
        RECT 4.400 562.000 1795.600 562.720 ;
        RECT 4.000 561.320 1795.600 562.000 ;
        RECT 4.000 509.680 1796.000 561.320 ;
        RECT 4.000 508.280 1795.600 509.680 ;
        RECT 4.000 487.920 1796.000 508.280 ;
        RECT 4.400 486.520 1796.000 487.920 ;
        RECT 4.000 455.960 1796.000 486.520 ;
        RECT 4.000 454.560 1795.600 455.960 ;
        RECT 4.000 413.120 1796.000 454.560 ;
        RECT 4.400 411.720 1796.000 413.120 ;
        RECT 4.000 402.240 1796.000 411.720 ;
        RECT 4.000 400.840 1795.600 402.240 ;
        RECT 4.000 348.520 1796.000 400.840 ;
        RECT 4.000 347.120 1795.600 348.520 ;
        RECT 4.000 338.320 1796.000 347.120 ;
        RECT 4.400 336.920 1796.000 338.320 ;
        RECT 4.000 294.800 1796.000 336.920 ;
        RECT 4.000 293.400 1795.600 294.800 ;
        RECT 4.000 262.840 1796.000 293.400 ;
        RECT 4.400 261.440 1796.000 262.840 ;
        RECT 4.000 241.760 1796.000 261.440 ;
        RECT 4.000 240.360 1795.600 241.760 ;
        RECT 4.000 188.040 1796.000 240.360 ;
        RECT 4.400 186.640 1795.600 188.040 ;
        RECT 4.000 134.320 1796.000 186.640 ;
        RECT 4.000 132.920 1795.600 134.320 ;
        RECT 4.000 113.240 1796.000 132.920 ;
        RECT 4.400 111.840 1796.000 113.240 ;
        RECT 4.000 80.600 1796.000 111.840 ;
        RECT 4.000 79.200 1795.600 80.600 ;
        RECT 4.000 38.440 1796.000 79.200 ;
        RECT 4.400 37.040 1796.000 38.440 ;
        RECT 4.000 27.560 1796.000 37.040 ;
        RECT 4.000 26.160 1795.600 27.560 ;
        RECT 4.000 10.715 1796.000 26.160 ;
      LAYER met4 ;
        RECT 25.135 11.735 97.440 1484.265 ;
        RECT 99.840 11.735 174.240 1484.265 ;
        RECT 176.640 11.735 251.040 1484.265 ;
        RECT 253.440 11.735 327.840 1484.265 ;
        RECT 330.240 11.735 404.640 1484.265 ;
        RECT 407.040 11.735 481.440 1484.265 ;
        RECT 483.840 11.735 558.240 1484.265 ;
        RECT 560.640 11.735 635.040 1484.265 ;
        RECT 637.440 11.735 711.840 1484.265 ;
        RECT 714.240 11.735 788.640 1484.265 ;
        RECT 791.040 11.735 865.440 1484.265 ;
        RECT 867.840 11.735 942.240 1484.265 ;
        RECT 944.640 11.735 1019.040 1484.265 ;
        RECT 1021.440 11.735 1095.840 1484.265 ;
        RECT 1098.240 11.735 1172.640 1484.265 ;
        RECT 1175.040 11.735 1249.440 1484.265 ;
        RECT 1251.840 11.735 1326.240 1484.265 ;
        RECT 1328.640 11.735 1403.040 1484.265 ;
        RECT 1405.440 11.735 1479.840 1484.265 ;
        RECT 1482.240 11.735 1556.640 1484.265 ;
        RECT 1559.040 11.735 1633.440 1484.265 ;
        RECT 1635.840 11.735 1710.240 1484.265 ;
        RECT 1712.640 11.735 1774.385 1484.265 ;
  END
END custom_sram
END LIBRARY

