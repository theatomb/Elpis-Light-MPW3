VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO custom_sram
  CLASS BLOCK ;
  FOREIGN custom_sram ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 1500.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 35.400 1800.000 36.000 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 0.000 956.250 4.000 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 1496.000 642.990 1500.000 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 606.600 1800.000 607.200 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 1496.000 814.570 1500.000 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 749.400 1800.000 750.000 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.160 4.000 924.760 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 4.000 975.080 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 4.000 1024.720 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 820.800 1800.000 821.400 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 178.200 1800.000 178.800 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 249.600 1800.000 250.200 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 1496.000 471.410 1500.000 ;
    END
  END a[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END clk
  PIN csb0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END csb0_to_sram
  PIN d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END d[0]
  PIN d[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END d[10]
  PIN d[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END d[11]
  PIN d[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 1496.000 728.550 1500.000 ;
    END
  END d[12]
  PIN d[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.200 4.000 824.800 ;
    END
  END d[13]
  PIN d[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 678.000 1800.000 678.600 ;
    END
  END d[14]
  PIN d[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END d[15]
  PIN d[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 0.000 1406.130 4.000 ;
    END
  END d[16]
  PIN d[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.550 0.000 1518.830 4.000 ;
    END
  END d[17]
  PIN d[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END d[18]
  PIN d[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 1496.000 1157.270 1500.000 ;
    END
  END d[19]
  PIN d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 1496.000 43.150 1500.000 ;
    END
  END d[1]
  PIN d[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1174.400 4.000 1175.000 ;
    END
  END d[20]
  PIN d[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.570 1496.000 1328.850 1500.000 ;
    END
  END d[21]
  PIN d[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.130 1496.000 1414.410 1500.000 ;
    END
  END d[22]
  PIN d[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.040 4.000 1224.640 ;
    END
  END d[23]
  PIN d[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1274.360 4.000 1274.960 ;
    END
  END d[24]
  PIN d[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 1496.000 1499.970 1500.000 ;
    END
  END d[25]
  PIN d[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.490 0.000 1743.770 4.000 ;
    END
  END d[26]
  PIN d[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1249.200 1800.000 1249.800 ;
    END
  END d[27]
  PIN d[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1324.000 4.000 1324.600 ;
    END
  END d[28]
  PIN d[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1392.000 1800.000 1392.600 ;
    END
  END d[29]
  PIN d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 1496.000 214.270 1500.000 ;
    END
  END d[2]
  PIN d[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1374.320 4.000 1374.920 ;
    END
  END d[30]
  PIN d[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1474.280 4.000 1474.880 ;
    END
  END d[31]
  PIN d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END d[3]
  PIN d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END d[4]
  PIN d[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END d[5]
  PIN d[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 1496.000 300.290 1500.000 ;
    END
  END d[6]
  PIN d[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 321.000 1800.000 321.600 ;
    END
  END d[7]
  PIN d[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 1496.000 385.850 1500.000 ;
    END
  END d[8]
  PIN d[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 1496.000 557.430 1500.000 ;
    END
  END d[9]
  PIN q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 106.800 1800.000 107.400 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 535.200 1800.000 535.800 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.670 0.000 1068.950 4.000 ;
    END
  END q[11]
  PIN q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 774.560 4.000 775.160 ;
    END
  END q[12]
  PIN q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 874.520 4.000 875.120 ;
    END
  END q[13]
  PIN q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1496.000 900.130 1500.000 ;
    END
  END q[14]
  PIN q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.610 0.000 1293.890 4.000 ;
    END
  END q[15]
  PIN q[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 1496.000 985.690 1500.000 ;
    END
  END q[16]
  PIN q[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 1496.000 1071.710 1500.000 ;
    END
  END q[17]
  PIN q[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.080 4.000 1124.680 ;
    END
  END q[18]
  PIN q[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 1496.000 1242.830 1500.000 ;
    END
  END q[19]
  PIN q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 1496.000 128.710 1500.000 ;
    END
  END q[1]
  PIN q[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 892.200 1800.000 892.800 ;
    END
  END q[20]
  PIN q[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 963.600 1800.000 964.200 ;
    END
  END q[21]
  PIN q[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1035.000 1800.000 1035.600 ;
    END
  END q[22]
  PIN q[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.790 0.000 1631.070 4.000 ;
    END
  END q[23]
  PIN q[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1106.400 1800.000 1107.000 ;
    END
  END q[24]
  PIN q[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.710 1496.000 1585.990 1500.000 ;
    END
  END q[25]
  PIN q[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1177.800 1800.000 1178.400 ;
    END
  END q[26]
  PIN q[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1320.600 1800.000 1321.200 ;
    END
  END q[27]
  PIN q[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 1496.000 1671.550 1500.000 ;
    END
  END q[28]
  PIN q[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.830 1496.000 1757.110 1500.000 ;
    END
  END q[29]
  PIN q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 4.000 325.000 ;
    END
  END q[2]
  PIN q[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1423.960 4.000 1424.560 ;
    END
  END q[30]
  PIN q[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1463.400 1800.000 1464.000 ;
    END
  END q[31]
  PIN q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 392.400 1800.000 393.000 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 463.800 1800.000 464.400 ;
    END
  END q[9]
  PIN spare_wen0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1488.080 ;
    END
  END vssd1
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END we
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1797.075 1487.925 ;
      LAYER met1 ;
        RECT 5.520 10.240 1797.135 1488.820 ;
      LAYER met2 ;
        RECT 6.600 1495.720 42.590 1496.410 ;
        RECT 43.430 1495.720 128.150 1496.410 ;
        RECT 128.990 1495.720 213.710 1496.410 ;
        RECT 214.550 1495.720 299.730 1496.410 ;
        RECT 300.570 1495.720 385.290 1496.410 ;
        RECT 386.130 1495.720 470.850 1496.410 ;
        RECT 471.690 1495.720 556.870 1496.410 ;
        RECT 557.710 1495.720 642.430 1496.410 ;
        RECT 643.270 1495.720 727.990 1496.410 ;
        RECT 728.830 1495.720 814.010 1496.410 ;
        RECT 814.850 1495.720 899.570 1496.410 ;
        RECT 900.410 1495.720 985.130 1496.410 ;
        RECT 985.970 1495.720 1071.150 1496.410 ;
        RECT 1071.990 1495.720 1156.710 1496.410 ;
        RECT 1157.550 1495.720 1242.270 1496.410 ;
        RECT 1243.110 1495.720 1328.290 1496.410 ;
        RECT 1329.130 1495.720 1413.850 1496.410 ;
        RECT 1414.690 1495.720 1499.410 1496.410 ;
        RECT 1500.250 1495.720 1585.430 1496.410 ;
        RECT 1586.270 1495.720 1670.990 1496.410 ;
        RECT 1671.830 1495.720 1756.550 1496.410 ;
        RECT 1757.390 1495.720 1795.290 1496.410 ;
        RECT 6.600 4.280 1795.290 1495.720 ;
        RECT 6.600 3.670 55.930 4.280 ;
        RECT 56.770 3.670 168.170 4.280 ;
        RECT 169.010 3.670 280.870 4.280 ;
        RECT 281.710 3.670 393.110 4.280 ;
        RECT 393.950 3.670 505.810 4.280 ;
        RECT 506.650 3.670 618.050 4.280 ;
        RECT 618.890 3.670 730.750 4.280 ;
        RECT 731.590 3.670 842.990 4.280 ;
        RECT 843.830 3.670 955.690 4.280 ;
        RECT 956.530 3.670 1068.390 4.280 ;
        RECT 1069.230 3.670 1180.630 4.280 ;
        RECT 1181.470 3.670 1293.330 4.280 ;
        RECT 1294.170 3.670 1405.570 4.280 ;
        RECT 1406.410 3.670 1518.270 4.280 ;
        RECT 1519.110 3.670 1630.510 4.280 ;
        RECT 1631.350 3.670 1743.210 4.280 ;
        RECT 1744.050 3.670 1795.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 1475.280 1796.000 1488.005 ;
        RECT 4.400 1473.880 1796.000 1475.280 ;
        RECT 4.000 1464.400 1796.000 1473.880 ;
        RECT 4.000 1463.000 1795.600 1464.400 ;
        RECT 4.000 1424.960 1796.000 1463.000 ;
        RECT 4.400 1423.560 1796.000 1424.960 ;
        RECT 4.000 1393.000 1796.000 1423.560 ;
        RECT 4.000 1391.600 1795.600 1393.000 ;
        RECT 4.000 1375.320 1796.000 1391.600 ;
        RECT 4.400 1373.920 1796.000 1375.320 ;
        RECT 4.000 1325.000 1796.000 1373.920 ;
        RECT 4.400 1323.600 1796.000 1325.000 ;
        RECT 4.000 1321.600 1796.000 1323.600 ;
        RECT 4.000 1320.200 1795.600 1321.600 ;
        RECT 4.000 1275.360 1796.000 1320.200 ;
        RECT 4.400 1273.960 1796.000 1275.360 ;
        RECT 4.000 1250.200 1796.000 1273.960 ;
        RECT 4.000 1248.800 1795.600 1250.200 ;
        RECT 4.000 1225.040 1796.000 1248.800 ;
        RECT 4.400 1223.640 1796.000 1225.040 ;
        RECT 4.000 1178.800 1796.000 1223.640 ;
        RECT 4.000 1177.400 1795.600 1178.800 ;
        RECT 4.000 1175.400 1796.000 1177.400 ;
        RECT 4.400 1174.000 1796.000 1175.400 ;
        RECT 4.000 1125.080 1796.000 1174.000 ;
        RECT 4.400 1123.680 1796.000 1125.080 ;
        RECT 4.000 1107.400 1796.000 1123.680 ;
        RECT 4.000 1106.000 1795.600 1107.400 ;
        RECT 4.000 1075.440 1796.000 1106.000 ;
        RECT 4.400 1074.040 1796.000 1075.440 ;
        RECT 4.000 1036.000 1796.000 1074.040 ;
        RECT 4.000 1034.600 1795.600 1036.000 ;
        RECT 4.000 1025.120 1796.000 1034.600 ;
        RECT 4.400 1023.720 1796.000 1025.120 ;
        RECT 4.000 975.480 1796.000 1023.720 ;
        RECT 4.400 974.080 1796.000 975.480 ;
        RECT 4.000 964.600 1796.000 974.080 ;
        RECT 4.000 963.200 1795.600 964.600 ;
        RECT 4.000 925.160 1796.000 963.200 ;
        RECT 4.400 923.760 1796.000 925.160 ;
        RECT 4.000 893.200 1796.000 923.760 ;
        RECT 4.000 891.800 1795.600 893.200 ;
        RECT 4.000 875.520 1796.000 891.800 ;
        RECT 4.400 874.120 1796.000 875.520 ;
        RECT 4.000 825.200 1796.000 874.120 ;
        RECT 4.400 823.800 1796.000 825.200 ;
        RECT 4.000 821.800 1796.000 823.800 ;
        RECT 4.000 820.400 1795.600 821.800 ;
        RECT 4.000 775.560 1796.000 820.400 ;
        RECT 4.400 774.160 1796.000 775.560 ;
        RECT 4.000 750.400 1796.000 774.160 ;
        RECT 4.000 749.000 1795.600 750.400 ;
        RECT 4.000 725.240 1796.000 749.000 ;
        RECT 4.400 723.840 1796.000 725.240 ;
        RECT 4.000 679.000 1796.000 723.840 ;
        RECT 4.000 677.600 1795.600 679.000 ;
        RECT 4.000 674.920 1796.000 677.600 ;
        RECT 4.400 673.520 1796.000 674.920 ;
        RECT 4.000 625.280 1796.000 673.520 ;
        RECT 4.400 623.880 1796.000 625.280 ;
        RECT 4.000 607.600 1796.000 623.880 ;
        RECT 4.000 606.200 1795.600 607.600 ;
        RECT 4.000 574.960 1796.000 606.200 ;
        RECT 4.400 573.560 1796.000 574.960 ;
        RECT 4.000 536.200 1796.000 573.560 ;
        RECT 4.000 534.800 1795.600 536.200 ;
        RECT 4.000 525.320 1796.000 534.800 ;
        RECT 4.400 523.920 1796.000 525.320 ;
        RECT 4.000 475.000 1796.000 523.920 ;
        RECT 4.400 473.600 1796.000 475.000 ;
        RECT 4.000 464.800 1796.000 473.600 ;
        RECT 4.000 463.400 1795.600 464.800 ;
        RECT 4.000 425.360 1796.000 463.400 ;
        RECT 4.400 423.960 1796.000 425.360 ;
        RECT 4.000 393.400 1796.000 423.960 ;
        RECT 4.000 392.000 1795.600 393.400 ;
        RECT 4.000 375.040 1796.000 392.000 ;
        RECT 4.400 373.640 1796.000 375.040 ;
        RECT 4.000 325.400 1796.000 373.640 ;
        RECT 4.400 324.000 1796.000 325.400 ;
        RECT 4.000 322.000 1796.000 324.000 ;
        RECT 4.000 320.600 1795.600 322.000 ;
        RECT 4.000 275.080 1796.000 320.600 ;
        RECT 4.400 273.680 1796.000 275.080 ;
        RECT 4.000 250.600 1796.000 273.680 ;
        RECT 4.000 249.200 1795.600 250.600 ;
        RECT 4.000 225.440 1796.000 249.200 ;
        RECT 4.400 224.040 1796.000 225.440 ;
        RECT 4.000 179.200 1796.000 224.040 ;
        RECT 4.000 177.800 1795.600 179.200 ;
        RECT 4.000 175.120 1796.000 177.800 ;
        RECT 4.400 173.720 1796.000 175.120 ;
        RECT 4.000 125.480 1796.000 173.720 ;
        RECT 4.400 124.080 1796.000 125.480 ;
        RECT 4.000 107.800 1796.000 124.080 ;
        RECT 4.000 106.400 1795.600 107.800 ;
        RECT 4.000 75.160 1796.000 106.400 ;
        RECT 4.400 73.760 1796.000 75.160 ;
        RECT 4.000 36.400 1796.000 73.760 ;
        RECT 4.000 35.000 1795.600 36.400 ;
        RECT 4.000 25.520 1796.000 35.000 ;
        RECT 4.400 24.120 1796.000 25.520 ;
        RECT 4.000 10.715 1796.000 24.120 ;
      LAYER met4 ;
        RECT 51.815 53.895 97.440 1486.305 ;
        RECT 99.840 53.895 174.240 1486.305 ;
        RECT 176.640 53.895 251.040 1486.305 ;
        RECT 253.440 53.895 327.840 1486.305 ;
        RECT 330.240 53.895 404.640 1486.305 ;
        RECT 407.040 53.895 481.440 1486.305 ;
        RECT 483.840 53.895 558.240 1486.305 ;
        RECT 560.640 53.895 635.040 1486.305 ;
        RECT 637.440 53.895 711.840 1486.305 ;
        RECT 714.240 53.895 788.640 1486.305 ;
        RECT 791.040 53.895 865.440 1486.305 ;
        RECT 867.840 53.895 942.240 1486.305 ;
        RECT 944.640 53.895 1019.040 1486.305 ;
        RECT 1021.440 53.895 1095.840 1486.305 ;
        RECT 1098.240 53.895 1172.640 1486.305 ;
        RECT 1175.040 53.895 1249.440 1486.305 ;
        RECT 1251.840 53.895 1326.240 1486.305 ;
        RECT 1328.640 53.895 1403.040 1486.305 ;
        RECT 1405.440 53.895 1479.840 1486.305 ;
        RECT 1482.240 53.895 1556.640 1486.305 ;
        RECT 1559.040 53.895 1633.440 1486.305 ;
        RECT 1635.840 53.895 1710.240 1486.305 ;
        RECT 1712.640 53.895 1786.345 1486.305 ;
  END
END custom_sram
END LIBRARY

