VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 1496.000 104.790 1500.000 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1317.880 4.000 1318.480 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.510 1496.000 1346.790 1500.000 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.930 0.000 1244.210 4.000 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1171.680 1500.000 1172.280 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1333.520 4.000 1334.120 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.160 4.000 1349.760 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.610 0.000 1293.890 4.000 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 0.000 1309.990 4.000 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1235.600 1500.000 1236.200 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.910 1496.000 1411.190 1500.000 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 199.960 1500.000 200.560 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.270 0.000 1326.550 4.000 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 0.000 1343.110 4.000 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.390 0.000 1359.670 4.000 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1277.760 1500.000 1278.360 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.610 0.000 1408.890 4.000 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 1496.000 1427.290 1500.000 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1319.920 1500.000 1320.520 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.110 1496.000 1443.390 1500.000 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1362.080 1500.000 1362.680 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.170 0.000 1425.450 4.000 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 1496.000 346.750 1500.000 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.730 0.000 1442.010 4.000 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1444.360 4.000 1444.960 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.210 1496.000 1459.490 1500.000 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1425.320 1500.000 1425.920 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1467.480 1500.000 1468.080 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1488.560 1500.000 1489.160 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 1496.000 1491.690 1500.000 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 221.040 1500.000 221.640 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 1496.000 508.210 1500.000 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 1496.000 540.410 1500.000 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 52.400 1500.000 53.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 1496.000 572.610 1500.000 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 1496.000 588.710 1500.000 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 432.520 1500.000 433.120 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 1496.000 620.910 1500.000 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 1496.000 653.110 1500.000 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 495.760 1500.000 496.360 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 516.840 1500.000 517.440 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 1496.000 701.410 1500.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 537.920 1500.000 538.520 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 1496.000 733.610 1500.000 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 559.000 1500.000 559.600 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 891.520 4.000 892.120 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 1496.000 169.190 1500.000 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 580.080 1500.000 580.680 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 1496.000 782.370 1500.000 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.160 4.000 907.760 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 601.160 1500.000 601.760 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.800 4.000 923.400 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 1496.000 798.470 1500.000 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 1496.000 846.770 1500.000 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 1496.000 878.970 1500.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.760 4.000 955.360 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 0.000 799.390 4.000 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 0.000 865.170 4.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 1496.000 927.270 1500.000 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 644.000 1500.000 644.600 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 1496.000 943.370 1500.000 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.680 4.000 1002.280 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.000 4.000 1018.600 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 94.560 1500.000 95.160 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 686.160 1500.000 686.760 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 1496.000 991.670 1500.000 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.950 1496.000 1008.230 1500.000 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 770.480 1500.000 771.080 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 791.560 1500.000 792.160 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1496.000 1040.430 1500.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.280 4.000 1049.880 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 833.720 1500.000 834.320 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 4.000 1065.520 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 1496.000 217.490 1500.000 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1496.000 1072.630 1500.000 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.550 1496.000 1104.830 1500.000 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 1496.000 1120.930 1500.000 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1112.520 4.000 1113.120 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 1496.000 1153.130 1500.000 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 1496.000 1169.230 1500.000 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 1496.000 1185.330 1500.000 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 1496.000 266.250 1500.000 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1128.160 4.000 1128.760 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1143.800 4.000 1144.400 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 918.720 1500.000 919.320 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1160.120 4.000 1160.720 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 939.800 1500.000 940.400 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 0.000 1112.190 4.000 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.350 1496.000 1233.630 1500.000 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 981.960 1500.000 982.560 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.040 4.000 1207.640 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.000 4.000 1239.600 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.590 0.000 1161.870 4.000 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1254.640 4.000 1255.240 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 0.000 1227.650 4.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.280 4.000 1270.880 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.110 1496.000 1282.390 1500.000 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1045.200 1500.000 1045.800 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.920 4.000 1286.520 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 1496.000 1314.590 1500.000 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1108.440 1500.000 1109.040 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 10.240 1500.000 10.840 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 1496.000 362.850 1500.000 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 1496.000 443.350 1500.000 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 263.200 1500.000 263.800 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 284.280 1500.000 284.880 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 528.400 4.000 529.000 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 1496.000 120.890 1500.000 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.880 4.000 655.480 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 1496.000 669.210 1500.000 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 4.000 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 1496.000 185.290 1500.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 115.640 1500.000 116.240 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 1496.000 298.450 1500.000 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 157.800 1500.000 158.400 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 1496.000 40.390 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 1496.000 88.690 1500.000 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 1496.000 72.590 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 1496.000 56.490 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 242.120 1500.000 242.720 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 1496.000 411.150 1500.000 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 305.360 1500.000 305.960 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 1496.000 556.510 1500.000 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 1496.000 136.990 1500.000 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 73.480 1500.000 74.080 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 1496.000 1330.690 1500.000 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1150.600 1500.000 1151.200 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.490 0.000 1260.770 4.000 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.610 1496.000 1362.890 1500.000 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.050 0.000 1277.330 4.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1192.760 1500.000 1193.360 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1214.520 1500.000 1215.120 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 1496.000 1378.990 1500.000 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.810 1496.000 1395.090 1500.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1365.480 4.000 1366.080 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1381.120 4.000 1381.720 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1256.680 1500.000 1257.280 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.950 0.000 1376.230 4.000 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.510 0.000 1392.790 4.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1298.840 1500.000 1299.440 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1396.760 4.000 1397.360 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1341.000 1500.000 1341.600 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1412.400 4.000 1413.000 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1383.160 1500.000 1383.760 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.040 4.000 1428.640 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1404.240 1500.000 1404.840 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.290 0.000 1458.570 4.000 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 1496.000 1475.590 1500.000 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1446.400 1500.000 1447.000 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1460.000 4.000 1460.600 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 0.000 1491.690 4.000 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1475.640 4.000 1476.240 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.280 4.000 1491.880 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 1496.000 395.050 1500.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 1496.000 427.250 1500.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 1496.000 459.450 1500.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 1496.000 475.550 1500.000 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 1496.000 524.310 1500.000 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 1496.000 153.090 1500.000 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 348.200 1500.000 348.800 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 369.280 1500.000 369.880 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1496.000 604.810 1500.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 453.600 1500.000 454.200 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 1496.000 637.010 1500.000 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 474.680 1500.000 475.280 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.760 4.000 734.360 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 1496.000 685.310 1500.000 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 1496.000 717.510 1500.000 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 0.000 683.930 4.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.920 4.000 844.520 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 1496.000 749.710 1500.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 1496.000 766.270 1500.000 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 622.920 1500.000 623.520 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 1496.000 814.570 1500.000 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 1496.000 830.670 1500.000 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 1496.000 862.870 1500.000 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 1496.000 895.070 1500.000 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 1496.000 911.170 1500.000 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 0.000 848.610 4.000 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 0.000 898.290 4.000 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 970.400 4.000 971.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 1496.000 959.470 1500.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 1496.000 975.570 1500.000 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 665.080 1500.000 665.680 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.110 0.000 914.390 4.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 707.240 1500.000 707.840 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 728.320 1500.000 728.920 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 749.400 1500.000 750.000 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 1496.000 1024.330 1500.000 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 812.640 1500.000 813.240 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 4.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 0.000 964.070 4.000 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 854.800 1500.000 855.400 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 1496.000 233.590 1500.000 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 1496.000 1056.530 1500.000 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.450 1496.000 1088.730 1500.000 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 0.000 997.190 4.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.880 4.000 1097.480 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 875.880 1500.000 876.480 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 1496.000 1137.030 1500.000 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 0.000 1079.530 4.000 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 0.000 1096.090 4.000 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 1496.000 1201.430 1500.000 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 896.960 1500.000 897.560 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.250 1496.000 1217.530 1500.000 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1175.760 4.000 1176.360 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1191.400 4.000 1192.000 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 0.000 1128.750 4.000 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 960.880 1500.000 961.480 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1003.040 1500.000 1003.640 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1223.360 4.000 1223.960 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.030 0.000 1145.310 4.000 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 1496.000 314.550 1500.000 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.150 0.000 1178.430 4.000 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 0.000 1194.990 4.000 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 1496.000 1249.730 1500.000 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1024.120 1500.000 1024.720 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 1496.000 1266.290 1500.000 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 1496.000 1298.490 1500.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1066.280 1500.000 1066.880 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1087.360 1500.000 1087.960 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.240 4.000 1302.840 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1129.520 1500.000 1130.120 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 178.880 1500.000 179.480 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 1496.000 8.190 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 1496.000 24.290 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 31.320 1500.000 31.920 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 1496.000 330.650 1500.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 1496.000 378.950 1500.000 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 1496.000 491.650 1500.000 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 327.120 1500.000 327.720 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 390.360 1500.000 390.960 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 411.440 1500.000 412.040 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 1496.000 201.390 1500.000 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 1496.000 249.690 1500.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 1496.000 282.350 1500.000 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 136.720 1500.000 137.320 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.080 1488.080 ;
      LAYER met2 ;
        RECT 6.990 1495.720 7.630 1496.410 ;
        RECT 8.470 1495.720 23.730 1496.410 ;
        RECT 24.570 1495.720 39.830 1496.410 ;
        RECT 40.670 1495.720 55.930 1496.410 ;
        RECT 56.770 1495.720 72.030 1496.410 ;
        RECT 72.870 1495.720 88.130 1496.410 ;
        RECT 88.970 1495.720 104.230 1496.410 ;
        RECT 105.070 1495.720 120.330 1496.410 ;
        RECT 121.170 1495.720 136.430 1496.410 ;
        RECT 137.270 1495.720 152.530 1496.410 ;
        RECT 153.370 1495.720 168.630 1496.410 ;
        RECT 169.470 1495.720 184.730 1496.410 ;
        RECT 185.570 1495.720 200.830 1496.410 ;
        RECT 201.670 1495.720 216.930 1496.410 ;
        RECT 217.770 1495.720 233.030 1496.410 ;
        RECT 233.870 1495.720 249.130 1496.410 ;
        RECT 249.970 1495.720 265.690 1496.410 ;
        RECT 266.530 1495.720 281.790 1496.410 ;
        RECT 282.630 1495.720 297.890 1496.410 ;
        RECT 298.730 1495.720 313.990 1496.410 ;
        RECT 314.830 1495.720 330.090 1496.410 ;
        RECT 330.930 1495.720 346.190 1496.410 ;
        RECT 347.030 1495.720 362.290 1496.410 ;
        RECT 363.130 1495.720 378.390 1496.410 ;
        RECT 379.230 1495.720 394.490 1496.410 ;
        RECT 395.330 1495.720 410.590 1496.410 ;
        RECT 411.430 1495.720 426.690 1496.410 ;
        RECT 427.530 1495.720 442.790 1496.410 ;
        RECT 443.630 1495.720 458.890 1496.410 ;
        RECT 459.730 1495.720 474.990 1496.410 ;
        RECT 475.830 1495.720 491.090 1496.410 ;
        RECT 491.930 1495.720 507.650 1496.410 ;
        RECT 508.490 1495.720 523.750 1496.410 ;
        RECT 524.590 1495.720 539.850 1496.410 ;
        RECT 540.690 1495.720 555.950 1496.410 ;
        RECT 556.790 1495.720 572.050 1496.410 ;
        RECT 572.890 1495.720 588.150 1496.410 ;
        RECT 588.990 1495.720 604.250 1496.410 ;
        RECT 605.090 1495.720 620.350 1496.410 ;
        RECT 621.190 1495.720 636.450 1496.410 ;
        RECT 637.290 1495.720 652.550 1496.410 ;
        RECT 653.390 1495.720 668.650 1496.410 ;
        RECT 669.490 1495.720 684.750 1496.410 ;
        RECT 685.590 1495.720 700.850 1496.410 ;
        RECT 701.690 1495.720 716.950 1496.410 ;
        RECT 717.790 1495.720 733.050 1496.410 ;
        RECT 733.890 1495.720 749.150 1496.410 ;
        RECT 749.990 1495.720 765.710 1496.410 ;
        RECT 766.550 1495.720 781.810 1496.410 ;
        RECT 782.650 1495.720 797.910 1496.410 ;
        RECT 798.750 1495.720 814.010 1496.410 ;
        RECT 814.850 1495.720 830.110 1496.410 ;
        RECT 830.950 1495.720 846.210 1496.410 ;
        RECT 847.050 1495.720 862.310 1496.410 ;
        RECT 863.150 1495.720 878.410 1496.410 ;
        RECT 879.250 1495.720 894.510 1496.410 ;
        RECT 895.350 1495.720 910.610 1496.410 ;
        RECT 911.450 1495.720 926.710 1496.410 ;
        RECT 927.550 1495.720 942.810 1496.410 ;
        RECT 943.650 1495.720 958.910 1496.410 ;
        RECT 959.750 1495.720 975.010 1496.410 ;
        RECT 975.850 1495.720 991.110 1496.410 ;
        RECT 991.950 1495.720 1007.670 1496.410 ;
        RECT 1008.510 1495.720 1023.770 1496.410 ;
        RECT 1024.610 1495.720 1039.870 1496.410 ;
        RECT 1040.710 1495.720 1055.970 1496.410 ;
        RECT 1056.810 1495.720 1072.070 1496.410 ;
        RECT 1072.910 1495.720 1088.170 1496.410 ;
        RECT 1089.010 1495.720 1104.270 1496.410 ;
        RECT 1105.110 1495.720 1120.370 1496.410 ;
        RECT 1121.210 1495.720 1136.470 1496.410 ;
        RECT 1137.310 1495.720 1152.570 1496.410 ;
        RECT 1153.410 1495.720 1168.670 1496.410 ;
        RECT 1169.510 1495.720 1184.770 1496.410 ;
        RECT 1185.610 1495.720 1200.870 1496.410 ;
        RECT 1201.710 1495.720 1216.970 1496.410 ;
        RECT 1217.810 1495.720 1233.070 1496.410 ;
        RECT 1233.910 1495.720 1249.170 1496.410 ;
        RECT 1250.010 1495.720 1265.730 1496.410 ;
        RECT 1266.570 1495.720 1281.830 1496.410 ;
        RECT 1282.670 1495.720 1297.930 1496.410 ;
        RECT 1298.770 1495.720 1314.030 1496.410 ;
        RECT 1314.870 1495.720 1330.130 1496.410 ;
        RECT 1330.970 1495.720 1346.230 1496.410 ;
        RECT 1347.070 1495.720 1362.330 1496.410 ;
        RECT 1363.170 1495.720 1378.430 1496.410 ;
        RECT 1379.270 1495.720 1394.530 1496.410 ;
        RECT 1395.370 1495.720 1410.630 1496.410 ;
        RECT 1411.470 1495.720 1426.730 1496.410 ;
        RECT 1427.570 1495.720 1442.830 1496.410 ;
        RECT 1443.670 1495.720 1458.930 1496.410 ;
        RECT 1459.770 1495.720 1475.030 1496.410 ;
        RECT 1475.870 1495.720 1491.130 1496.410 ;
        RECT 6.990 4.280 1491.680 1495.720 ;
        RECT 6.990 4.000 7.630 4.280 ;
        RECT 8.470 4.000 23.730 4.280 ;
        RECT 24.570 4.000 40.290 4.280 ;
        RECT 41.130 4.000 56.850 4.280 ;
        RECT 57.690 4.000 73.410 4.280 ;
        RECT 74.250 4.000 89.970 4.280 ;
        RECT 90.810 4.000 106.530 4.280 ;
        RECT 107.370 4.000 122.630 4.280 ;
        RECT 123.470 4.000 139.190 4.280 ;
        RECT 140.030 4.000 155.750 4.280 ;
        RECT 156.590 4.000 172.310 4.280 ;
        RECT 173.150 4.000 188.870 4.280 ;
        RECT 189.710 4.000 205.430 4.280 ;
        RECT 206.270 4.000 221.530 4.280 ;
        RECT 222.370 4.000 238.090 4.280 ;
        RECT 238.930 4.000 254.650 4.280 ;
        RECT 255.490 4.000 271.210 4.280 ;
        RECT 272.050 4.000 287.770 4.280 ;
        RECT 288.610 4.000 304.330 4.280 ;
        RECT 305.170 4.000 320.430 4.280 ;
        RECT 321.270 4.000 336.990 4.280 ;
        RECT 337.830 4.000 353.550 4.280 ;
        RECT 354.390 4.000 370.110 4.280 ;
        RECT 370.950 4.000 386.670 4.280 ;
        RECT 387.510 4.000 403.230 4.280 ;
        RECT 404.070 4.000 419.330 4.280 ;
        RECT 420.170 4.000 435.890 4.280 ;
        RECT 436.730 4.000 452.450 4.280 ;
        RECT 453.290 4.000 469.010 4.280 ;
        RECT 469.850 4.000 485.570 4.280 ;
        RECT 486.410 4.000 502.130 4.280 ;
        RECT 502.970 4.000 518.230 4.280 ;
        RECT 519.070 4.000 534.790 4.280 ;
        RECT 535.630 4.000 551.350 4.280 ;
        RECT 552.190 4.000 567.910 4.280 ;
        RECT 568.750 4.000 584.470 4.280 ;
        RECT 585.310 4.000 601.030 4.280 ;
        RECT 601.870 4.000 617.130 4.280 ;
        RECT 617.970 4.000 633.690 4.280 ;
        RECT 634.530 4.000 650.250 4.280 ;
        RECT 651.090 4.000 666.810 4.280 ;
        RECT 667.650 4.000 683.370 4.280 ;
        RECT 684.210 4.000 699.930 4.280 ;
        RECT 700.770 4.000 716.030 4.280 ;
        RECT 716.870 4.000 732.590 4.280 ;
        RECT 733.430 4.000 749.150 4.280 ;
        RECT 749.990 4.000 765.710 4.280 ;
        RECT 766.550 4.000 782.270 4.280 ;
        RECT 783.110 4.000 798.830 4.280 ;
        RECT 799.670 4.000 814.930 4.280 ;
        RECT 815.770 4.000 831.490 4.280 ;
        RECT 832.330 4.000 848.050 4.280 ;
        RECT 848.890 4.000 864.610 4.280 ;
        RECT 865.450 4.000 881.170 4.280 ;
        RECT 882.010 4.000 897.730 4.280 ;
        RECT 898.570 4.000 913.830 4.280 ;
        RECT 914.670 4.000 930.390 4.280 ;
        RECT 931.230 4.000 946.950 4.280 ;
        RECT 947.790 4.000 963.510 4.280 ;
        RECT 964.350 4.000 980.070 4.280 ;
        RECT 980.910 4.000 996.630 4.280 ;
        RECT 997.470 4.000 1012.730 4.280 ;
        RECT 1013.570 4.000 1029.290 4.280 ;
        RECT 1030.130 4.000 1045.850 4.280 ;
        RECT 1046.690 4.000 1062.410 4.280 ;
        RECT 1063.250 4.000 1078.970 4.280 ;
        RECT 1079.810 4.000 1095.530 4.280 ;
        RECT 1096.370 4.000 1111.630 4.280 ;
        RECT 1112.470 4.000 1128.190 4.280 ;
        RECT 1129.030 4.000 1144.750 4.280 ;
        RECT 1145.590 4.000 1161.310 4.280 ;
        RECT 1162.150 4.000 1177.870 4.280 ;
        RECT 1178.710 4.000 1194.430 4.280 ;
        RECT 1195.270 4.000 1210.530 4.280 ;
        RECT 1211.370 4.000 1227.090 4.280 ;
        RECT 1227.930 4.000 1243.650 4.280 ;
        RECT 1244.490 4.000 1260.210 4.280 ;
        RECT 1261.050 4.000 1276.770 4.280 ;
        RECT 1277.610 4.000 1293.330 4.280 ;
        RECT 1294.170 4.000 1309.430 4.280 ;
        RECT 1310.270 4.000 1325.990 4.280 ;
        RECT 1326.830 4.000 1342.550 4.280 ;
        RECT 1343.390 4.000 1359.110 4.280 ;
        RECT 1359.950 4.000 1375.670 4.280 ;
        RECT 1376.510 4.000 1392.230 4.280 ;
        RECT 1393.070 4.000 1408.330 4.280 ;
        RECT 1409.170 4.000 1424.890 4.280 ;
        RECT 1425.730 4.000 1441.450 4.280 ;
        RECT 1442.290 4.000 1458.010 4.280 ;
        RECT 1458.850 4.000 1474.570 4.280 ;
        RECT 1475.410 4.000 1491.130 4.280 ;
      LAYER met3 ;
        RECT 4.400 1490.880 1496.000 1491.745 ;
        RECT 4.000 1489.560 1496.000 1490.880 ;
        RECT 4.000 1488.160 1495.600 1489.560 ;
        RECT 4.000 1476.640 1496.000 1488.160 ;
        RECT 4.400 1475.240 1496.000 1476.640 ;
        RECT 4.000 1468.480 1496.000 1475.240 ;
        RECT 4.000 1467.080 1495.600 1468.480 ;
        RECT 4.000 1461.000 1496.000 1467.080 ;
        RECT 4.400 1459.600 1496.000 1461.000 ;
        RECT 4.000 1447.400 1496.000 1459.600 ;
        RECT 4.000 1446.000 1495.600 1447.400 ;
        RECT 4.000 1445.360 1496.000 1446.000 ;
        RECT 4.400 1443.960 1496.000 1445.360 ;
        RECT 4.000 1429.040 1496.000 1443.960 ;
        RECT 4.400 1427.640 1496.000 1429.040 ;
        RECT 4.000 1426.320 1496.000 1427.640 ;
        RECT 4.000 1424.920 1495.600 1426.320 ;
        RECT 4.000 1413.400 1496.000 1424.920 ;
        RECT 4.400 1412.000 1496.000 1413.400 ;
        RECT 4.000 1405.240 1496.000 1412.000 ;
        RECT 4.000 1403.840 1495.600 1405.240 ;
        RECT 4.000 1397.760 1496.000 1403.840 ;
        RECT 4.400 1396.360 1496.000 1397.760 ;
        RECT 4.000 1384.160 1496.000 1396.360 ;
        RECT 4.000 1382.760 1495.600 1384.160 ;
        RECT 4.000 1382.120 1496.000 1382.760 ;
        RECT 4.400 1380.720 1496.000 1382.120 ;
        RECT 4.000 1366.480 1496.000 1380.720 ;
        RECT 4.400 1365.080 1496.000 1366.480 ;
        RECT 4.000 1363.080 1496.000 1365.080 ;
        RECT 4.000 1361.680 1495.600 1363.080 ;
        RECT 4.000 1350.160 1496.000 1361.680 ;
        RECT 4.400 1348.760 1496.000 1350.160 ;
        RECT 4.000 1342.000 1496.000 1348.760 ;
        RECT 4.000 1340.600 1495.600 1342.000 ;
        RECT 4.000 1334.520 1496.000 1340.600 ;
        RECT 4.400 1333.120 1496.000 1334.520 ;
        RECT 4.000 1320.920 1496.000 1333.120 ;
        RECT 4.000 1319.520 1495.600 1320.920 ;
        RECT 4.000 1318.880 1496.000 1319.520 ;
        RECT 4.400 1317.480 1496.000 1318.880 ;
        RECT 4.000 1303.240 1496.000 1317.480 ;
        RECT 4.400 1301.840 1496.000 1303.240 ;
        RECT 4.000 1299.840 1496.000 1301.840 ;
        RECT 4.000 1298.440 1495.600 1299.840 ;
        RECT 4.000 1286.920 1496.000 1298.440 ;
        RECT 4.400 1285.520 1496.000 1286.920 ;
        RECT 4.000 1278.760 1496.000 1285.520 ;
        RECT 4.000 1277.360 1495.600 1278.760 ;
        RECT 4.000 1271.280 1496.000 1277.360 ;
        RECT 4.400 1269.880 1496.000 1271.280 ;
        RECT 4.000 1257.680 1496.000 1269.880 ;
        RECT 4.000 1256.280 1495.600 1257.680 ;
        RECT 4.000 1255.640 1496.000 1256.280 ;
        RECT 4.400 1254.240 1496.000 1255.640 ;
        RECT 4.000 1240.000 1496.000 1254.240 ;
        RECT 4.400 1238.600 1496.000 1240.000 ;
        RECT 4.000 1236.600 1496.000 1238.600 ;
        RECT 4.000 1235.200 1495.600 1236.600 ;
        RECT 4.000 1224.360 1496.000 1235.200 ;
        RECT 4.400 1222.960 1496.000 1224.360 ;
        RECT 4.000 1215.520 1496.000 1222.960 ;
        RECT 4.000 1214.120 1495.600 1215.520 ;
        RECT 4.000 1208.040 1496.000 1214.120 ;
        RECT 4.400 1206.640 1496.000 1208.040 ;
        RECT 4.000 1193.760 1496.000 1206.640 ;
        RECT 4.000 1192.400 1495.600 1193.760 ;
        RECT 4.400 1192.360 1495.600 1192.400 ;
        RECT 4.400 1191.000 1496.000 1192.360 ;
        RECT 4.000 1176.760 1496.000 1191.000 ;
        RECT 4.400 1175.360 1496.000 1176.760 ;
        RECT 4.000 1172.680 1496.000 1175.360 ;
        RECT 4.000 1171.280 1495.600 1172.680 ;
        RECT 4.000 1161.120 1496.000 1171.280 ;
        RECT 4.400 1159.720 1496.000 1161.120 ;
        RECT 4.000 1151.600 1496.000 1159.720 ;
        RECT 4.000 1150.200 1495.600 1151.600 ;
        RECT 4.000 1144.800 1496.000 1150.200 ;
        RECT 4.400 1143.400 1496.000 1144.800 ;
        RECT 4.000 1130.520 1496.000 1143.400 ;
        RECT 4.000 1129.160 1495.600 1130.520 ;
        RECT 4.400 1129.120 1495.600 1129.160 ;
        RECT 4.400 1127.760 1496.000 1129.120 ;
        RECT 4.000 1113.520 1496.000 1127.760 ;
        RECT 4.400 1112.120 1496.000 1113.520 ;
        RECT 4.000 1109.440 1496.000 1112.120 ;
        RECT 4.000 1108.040 1495.600 1109.440 ;
        RECT 4.000 1097.880 1496.000 1108.040 ;
        RECT 4.400 1096.480 1496.000 1097.880 ;
        RECT 4.000 1088.360 1496.000 1096.480 ;
        RECT 4.000 1086.960 1495.600 1088.360 ;
        RECT 4.000 1082.240 1496.000 1086.960 ;
        RECT 4.400 1080.840 1496.000 1082.240 ;
        RECT 4.000 1067.280 1496.000 1080.840 ;
        RECT 4.000 1065.920 1495.600 1067.280 ;
        RECT 4.400 1065.880 1495.600 1065.920 ;
        RECT 4.400 1064.520 1496.000 1065.880 ;
        RECT 4.000 1050.280 1496.000 1064.520 ;
        RECT 4.400 1048.880 1496.000 1050.280 ;
        RECT 4.000 1046.200 1496.000 1048.880 ;
        RECT 4.000 1044.800 1495.600 1046.200 ;
        RECT 4.000 1034.640 1496.000 1044.800 ;
        RECT 4.400 1033.240 1496.000 1034.640 ;
        RECT 4.000 1025.120 1496.000 1033.240 ;
        RECT 4.000 1023.720 1495.600 1025.120 ;
        RECT 4.000 1019.000 1496.000 1023.720 ;
        RECT 4.400 1017.600 1496.000 1019.000 ;
        RECT 4.000 1004.040 1496.000 1017.600 ;
        RECT 4.000 1002.680 1495.600 1004.040 ;
        RECT 4.400 1002.640 1495.600 1002.680 ;
        RECT 4.400 1001.280 1496.000 1002.640 ;
        RECT 4.000 987.040 1496.000 1001.280 ;
        RECT 4.400 985.640 1496.000 987.040 ;
        RECT 4.000 982.960 1496.000 985.640 ;
        RECT 4.000 981.560 1495.600 982.960 ;
        RECT 4.000 971.400 1496.000 981.560 ;
        RECT 4.400 970.000 1496.000 971.400 ;
        RECT 4.000 961.880 1496.000 970.000 ;
        RECT 4.000 960.480 1495.600 961.880 ;
        RECT 4.000 955.760 1496.000 960.480 ;
        RECT 4.400 954.360 1496.000 955.760 ;
        RECT 4.000 940.800 1496.000 954.360 ;
        RECT 4.000 940.120 1495.600 940.800 ;
        RECT 4.400 939.400 1495.600 940.120 ;
        RECT 4.400 938.720 1496.000 939.400 ;
        RECT 4.000 923.800 1496.000 938.720 ;
        RECT 4.400 922.400 1496.000 923.800 ;
        RECT 4.000 919.720 1496.000 922.400 ;
        RECT 4.000 918.320 1495.600 919.720 ;
        RECT 4.000 908.160 1496.000 918.320 ;
        RECT 4.400 906.760 1496.000 908.160 ;
        RECT 4.000 897.960 1496.000 906.760 ;
        RECT 4.000 896.560 1495.600 897.960 ;
        RECT 4.000 892.520 1496.000 896.560 ;
        RECT 4.400 891.120 1496.000 892.520 ;
        RECT 4.000 876.880 1496.000 891.120 ;
        RECT 4.400 875.480 1495.600 876.880 ;
        RECT 4.000 860.560 1496.000 875.480 ;
        RECT 4.400 859.160 1496.000 860.560 ;
        RECT 4.000 855.800 1496.000 859.160 ;
        RECT 4.000 854.400 1495.600 855.800 ;
        RECT 4.000 844.920 1496.000 854.400 ;
        RECT 4.400 843.520 1496.000 844.920 ;
        RECT 4.000 834.720 1496.000 843.520 ;
        RECT 4.000 833.320 1495.600 834.720 ;
        RECT 4.000 829.280 1496.000 833.320 ;
        RECT 4.400 827.880 1496.000 829.280 ;
        RECT 4.000 813.640 1496.000 827.880 ;
        RECT 4.400 812.240 1495.600 813.640 ;
        RECT 4.000 798.000 1496.000 812.240 ;
        RECT 4.400 796.600 1496.000 798.000 ;
        RECT 4.000 792.560 1496.000 796.600 ;
        RECT 4.000 791.160 1495.600 792.560 ;
        RECT 4.000 781.680 1496.000 791.160 ;
        RECT 4.400 780.280 1496.000 781.680 ;
        RECT 4.000 771.480 1496.000 780.280 ;
        RECT 4.000 770.080 1495.600 771.480 ;
        RECT 4.000 766.040 1496.000 770.080 ;
        RECT 4.400 764.640 1496.000 766.040 ;
        RECT 4.000 750.400 1496.000 764.640 ;
        RECT 4.400 749.000 1495.600 750.400 ;
        RECT 4.000 734.760 1496.000 749.000 ;
        RECT 4.400 733.360 1496.000 734.760 ;
        RECT 4.000 729.320 1496.000 733.360 ;
        RECT 4.000 727.920 1495.600 729.320 ;
        RECT 4.000 718.440 1496.000 727.920 ;
        RECT 4.400 717.040 1496.000 718.440 ;
        RECT 4.000 708.240 1496.000 717.040 ;
        RECT 4.000 706.840 1495.600 708.240 ;
        RECT 4.000 702.800 1496.000 706.840 ;
        RECT 4.400 701.400 1496.000 702.800 ;
        RECT 4.000 687.160 1496.000 701.400 ;
        RECT 4.400 685.760 1495.600 687.160 ;
        RECT 4.000 671.520 1496.000 685.760 ;
        RECT 4.400 670.120 1496.000 671.520 ;
        RECT 4.000 666.080 1496.000 670.120 ;
        RECT 4.000 664.680 1495.600 666.080 ;
        RECT 4.000 655.880 1496.000 664.680 ;
        RECT 4.400 654.480 1496.000 655.880 ;
        RECT 4.000 645.000 1496.000 654.480 ;
        RECT 4.000 643.600 1495.600 645.000 ;
        RECT 4.000 639.560 1496.000 643.600 ;
        RECT 4.400 638.160 1496.000 639.560 ;
        RECT 4.000 623.920 1496.000 638.160 ;
        RECT 4.400 622.520 1495.600 623.920 ;
        RECT 4.000 608.280 1496.000 622.520 ;
        RECT 4.400 606.880 1496.000 608.280 ;
        RECT 4.000 602.160 1496.000 606.880 ;
        RECT 4.000 600.760 1495.600 602.160 ;
        RECT 4.000 592.640 1496.000 600.760 ;
        RECT 4.400 591.240 1496.000 592.640 ;
        RECT 4.000 581.080 1496.000 591.240 ;
        RECT 4.000 579.680 1495.600 581.080 ;
        RECT 4.000 576.320 1496.000 579.680 ;
        RECT 4.400 574.920 1496.000 576.320 ;
        RECT 4.000 560.680 1496.000 574.920 ;
        RECT 4.400 560.000 1496.000 560.680 ;
        RECT 4.400 559.280 1495.600 560.000 ;
        RECT 4.000 558.600 1495.600 559.280 ;
        RECT 4.000 545.040 1496.000 558.600 ;
        RECT 4.400 543.640 1496.000 545.040 ;
        RECT 4.000 538.920 1496.000 543.640 ;
        RECT 4.000 537.520 1495.600 538.920 ;
        RECT 4.000 529.400 1496.000 537.520 ;
        RECT 4.400 528.000 1496.000 529.400 ;
        RECT 4.000 517.840 1496.000 528.000 ;
        RECT 4.000 516.440 1495.600 517.840 ;
        RECT 4.000 513.760 1496.000 516.440 ;
        RECT 4.400 512.360 1496.000 513.760 ;
        RECT 4.000 497.440 1496.000 512.360 ;
        RECT 4.400 496.760 1496.000 497.440 ;
        RECT 4.400 496.040 1495.600 496.760 ;
        RECT 4.000 495.360 1495.600 496.040 ;
        RECT 4.000 481.800 1496.000 495.360 ;
        RECT 4.400 480.400 1496.000 481.800 ;
        RECT 4.000 475.680 1496.000 480.400 ;
        RECT 4.000 474.280 1495.600 475.680 ;
        RECT 4.000 466.160 1496.000 474.280 ;
        RECT 4.400 464.760 1496.000 466.160 ;
        RECT 4.000 454.600 1496.000 464.760 ;
        RECT 4.000 453.200 1495.600 454.600 ;
        RECT 4.000 450.520 1496.000 453.200 ;
        RECT 4.400 449.120 1496.000 450.520 ;
        RECT 4.000 434.200 1496.000 449.120 ;
        RECT 4.400 433.520 1496.000 434.200 ;
        RECT 4.400 432.800 1495.600 433.520 ;
        RECT 4.000 432.120 1495.600 432.800 ;
        RECT 4.000 418.560 1496.000 432.120 ;
        RECT 4.400 417.160 1496.000 418.560 ;
        RECT 4.000 412.440 1496.000 417.160 ;
        RECT 4.000 411.040 1495.600 412.440 ;
        RECT 4.000 402.920 1496.000 411.040 ;
        RECT 4.400 401.520 1496.000 402.920 ;
        RECT 4.000 391.360 1496.000 401.520 ;
        RECT 4.000 389.960 1495.600 391.360 ;
        RECT 4.000 387.280 1496.000 389.960 ;
        RECT 4.400 385.880 1496.000 387.280 ;
        RECT 4.000 371.640 1496.000 385.880 ;
        RECT 4.400 370.280 1496.000 371.640 ;
        RECT 4.400 370.240 1495.600 370.280 ;
        RECT 4.000 368.880 1495.600 370.240 ;
        RECT 4.000 355.320 1496.000 368.880 ;
        RECT 4.400 353.920 1496.000 355.320 ;
        RECT 4.000 349.200 1496.000 353.920 ;
        RECT 4.000 347.800 1495.600 349.200 ;
        RECT 4.000 339.680 1496.000 347.800 ;
        RECT 4.400 338.280 1496.000 339.680 ;
        RECT 4.000 328.120 1496.000 338.280 ;
        RECT 4.000 326.720 1495.600 328.120 ;
        RECT 4.000 324.040 1496.000 326.720 ;
        RECT 4.400 322.640 1496.000 324.040 ;
        RECT 4.000 308.400 1496.000 322.640 ;
        RECT 4.400 307.000 1496.000 308.400 ;
        RECT 4.000 306.360 1496.000 307.000 ;
        RECT 4.000 304.960 1495.600 306.360 ;
        RECT 4.000 292.080 1496.000 304.960 ;
        RECT 4.400 290.680 1496.000 292.080 ;
        RECT 4.000 285.280 1496.000 290.680 ;
        RECT 4.000 283.880 1495.600 285.280 ;
        RECT 4.000 276.440 1496.000 283.880 ;
        RECT 4.400 275.040 1496.000 276.440 ;
        RECT 4.000 264.200 1496.000 275.040 ;
        RECT 4.000 262.800 1495.600 264.200 ;
        RECT 4.000 260.800 1496.000 262.800 ;
        RECT 4.400 259.400 1496.000 260.800 ;
        RECT 4.000 245.160 1496.000 259.400 ;
        RECT 4.400 243.760 1496.000 245.160 ;
        RECT 4.000 243.120 1496.000 243.760 ;
        RECT 4.000 241.720 1495.600 243.120 ;
        RECT 4.000 229.520 1496.000 241.720 ;
        RECT 4.400 228.120 1496.000 229.520 ;
        RECT 4.000 222.040 1496.000 228.120 ;
        RECT 4.000 220.640 1495.600 222.040 ;
        RECT 4.000 213.200 1496.000 220.640 ;
        RECT 4.400 211.800 1496.000 213.200 ;
        RECT 4.000 200.960 1496.000 211.800 ;
        RECT 4.000 199.560 1495.600 200.960 ;
        RECT 4.000 197.560 1496.000 199.560 ;
        RECT 4.400 196.160 1496.000 197.560 ;
        RECT 4.000 181.920 1496.000 196.160 ;
        RECT 4.400 180.520 1496.000 181.920 ;
        RECT 4.000 179.880 1496.000 180.520 ;
        RECT 4.000 178.480 1495.600 179.880 ;
        RECT 4.000 166.280 1496.000 178.480 ;
        RECT 4.400 164.880 1496.000 166.280 ;
        RECT 4.000 158.800 1496.000 164.880 ;
        RECT 4.000 157.400 1495.600 158.800 ;
        RECT 4.000 149.960 1496.000 157.400 ;
        RECT 4.400 148.560 1496.000 149.960 ;
        RECT 4.000 137.720 1496.000 148.560 ;
        RECT 4.000 136.320 1495.600 137.720 ;
        RECT 4.000 134.320 1496.000 136.320 ;
        RECT 4.400 132.920 1496.000 134.320 ;
        RECT 4.000 118.680 1496.000 132.920 ;
        RECT 4.400 117.280 1496.000 118.680 ;
        RECT 4.000 116.640 1496.000 117.280 ;
        RECT 4.000 115.240 1495.600 116.640 ;
        RECT 4.000 103.040 1496.000 115.240 ;
        RECT 4.400 101.640 1496.000 103.040 ;
        RECT 4.000 95.560 1496.000 101.640 ;
        RECT 4.000 94.160 1495.600 95.560 ;
        RECT 4.000 87.400 1496.000 94.160 ;
        RECT 4.400 86.000 1496.000 87.400 ;
        RECT 4.000 74.480 1496.000 86.000 ;
        RECT 4.000 73.080 1495.600 74.480 ;
        RECT 4.000 71.080 1496.000 73.080 ;
        RECT 4.400 69.680 1496.000 71.080 ;
        RECT 4.000 55.440 1496.000 69.680 ;
        RECT 4.400 54.040 1496.000 55.440 ;
        RECT 4.000 53.400 1496.000 54.040 ;
        RECT 4.000 52.000 1495.600 53.400 ;
        RECT 4.000 39.800 1496.000 52.000 ;
        RECT 4.400 38.400 1496.000 39.800 ;
        RECT 4.000 32.320 1496.000 38.400 ;
        RECT 4.000 30.920 1495.600 32.320 ;
        RECT 4.000 24.160 1496.000 30.920 ;
        RECT 4.400 22.760 1496.000 24.160 ;
        RECT 4.000 11.240 1496.000 22.760 ;
        RECT 4.000 9.840 1495.600 11.240 ;
        RECT 4.000 8.520 1496.000 9.840 ;
        RECT 4.400 7.655 1496.000 8.520 ;
      LAYER met4 ;
        RECT 58.255 11.055 97.440 1484.265 ;
        RECT 99.840 11.055 174.240 1484.265 ;
        RECT 176.640 11.055 251.040 1484.265 ;
        RECT 253.440 11.055 327.840 1484.265 ;
        RECT 330.240 11.055 404.640 1484.265 ;
        RECT 407.040 11.055 481.440 1484.265 ;
        RECT 483.840 11.055 558.240 1484.265 ;
        RECT 560.640 11.055 635.040 1484.265 ;
        RECT 637.440 11.055 711.840 1484.265 ;
        RECT 714.240 11.055 788.640 1484.265 ;
        RECT 791.040 11.055 865.440 1484.265 ;
        RECT 867.840 11.055 942.240 1484.265 ;
        RECT 944.640 11.055 1019.040 1484.265 ;
        RECT 1021.440 11.055 1064.145 1484.265 ;
  END
END core
END LIBRARY

