VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_controller
  CLASS BLOCK ;
  FOREIGN chip_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN addr0_to_sram[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END addr0_to_sram[0]
  PIN addr0_to_sram[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END addr0_to_sram[10]
  PIN addr0_to_sram[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END addr0_to_sram[11]
  PIN addr0_to_sram[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 396.000 71.670 400.000 ;
    END
  END addr0_to_sram[12]
  PIN addr0_to_sram[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 86.400 400.000 87.000 ;
    END
  END addr0_to_sram[13]
  PIN addr0_to_sram[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 396.000 87.770 400.000 ;
    END
  END addr0_to_sram[14]
  PIN addr0_to_sram[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END addr0_to_sram[15]
  PIN addr0_to_sram[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END addr0_to_sram[16]
  PIN addr0_to_sram[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END addr0_to_sram[17]
  PIN addr0_to_sram[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END addr0_to_sram[18]
  PIN addr0_to_sram[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 128.560 400.000 129.160 ;
    END
  END addr0_to_sram[19]
  PIN addr0_to_sram[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END addr0_to_sram[1]
  PIN addr0_to_sram[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 396.000 16.930 400.000 ;
    END
  END addr0_to_sram[2]
  PIN addr0_to_sram[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END addr0_to_sram[3]
  PIN addr0_to_sram[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 25.880 400.000 26.480 ;
    END
  END addr0_to_sram[4]
  PIN addr0_to_sram[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 396.000 37.630 400.000 ;
    END
  END addr0_to_sram[5]
  PIN addr0_to_sram[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 36.760 400.000 37.360 ;
    END
  END addr0_to_sram[6]
  PIN addr0_to_sram[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 42.880 400.000 43.480 ;
    END
  END addr0_to_sram[7]
  PIN addr0_to_sram[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 46.280 400.000 46.880 ;
    END
  END addr0_to_sram[8]
  PIN addr0_to_sram[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 57.160 400.000 57.760 ;
    END
  END addr0_to_sram[9]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 396.000 0.830 400.000 ;
    END
  END addr_in[0]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 72.120 400.000 72.720 ;
    END
  END addr_in[11]
  PIN addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 396.000 73.050 400.000 ;
    END
  END addr_in[12]
  PIN addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END addr_in[13]
  PIN addr_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END addr_in[14]
  PIN addr_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 396.000 92.370 400.000 ;
    END
  END addr_in[15]
  PIN addr_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END addr_in[16]
  PIN addr_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END addr_in[17]
  PIN addr_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 396.000 107.090 400.000 ;
    END
  END addr_in[18]
  PIN addr_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 396.000 115.370 400.000 ;
    END
  END addr_in[19]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 15.000 400.000 15.600 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 396.000 26.590 400.000 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 48.320 400.000 48.920 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END addr_in[9]
  PIN addr_to_core_mem[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END addr_to_core_mem[0]
  PIN addr_to_core_mem[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 396.000 65.230 400.000 ;
    END
  END addr_to_core_mem[10]
  PIN addr_to_core_mem[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END addr_to_core_mem[11]
  PIN addr_to_core_mem[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 396.000 74.890 400.000 ;
    END
  END addr_to_core_mem[12]
  PIN addr_to_core_mem[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 88.440 400.000 89.040 ;
    END
  END addr_to_core_mem[13]
  PIN addr_to_core_mem[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END addr_to_core_mem[14]
  PIN addr_to_core_mem[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END addr_to_core_mem[15]
  PIN addr_to_core_mem[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END addr_to_core_mem[16]
  PIN addr_to_core_mem[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END addr_to_core_mem[17]
  PIN addr_to_core_mem[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END addr_to_core_mem[18]
  PIN addr_to_core_mem[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END addr_to_core_mem[19]
  PIN addr_to_core_mem[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 9.560 400.000 10.160 ;
    END
  END addr_to_core_mem[1]
  PIN addr_to_core_mem[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END addr_to_core_mem[2]
  PIN addr_to_core_mem[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END addr_to_core_mem[3]
  PIN addr_to_core_mem[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END addr_to_core_mem[4]
  PIN addr_to_core_mem[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END addr_to_core_mem[5]
  PIN addr_to_core_mem[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 38.800 400.000 39.400 ;
    END
  END addr_to_core_mem[6]
  PIN addr_to_core_mem[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END addr_to_core_mem[7]
  PIN addr_to_core_mem[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END addr_to_core_mem[8]
  PIN addr_to_core_mem[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 396.000 63.390 400.000 ;
    END
  END addr_to_core_mem[9]
  PIN clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END clk
  PIN core0_data_print[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END core0_data_print[0]
  PIN core0_data_print[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END core0_data_print[10]
  PIN core0_data_print[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END core0_data_print[11]
  PIN core0_data_print[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 80.960 400.000 81.560 ;
    END
  END core0_data_print[12]
  PIN core0_data_print[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 90.480 400.000 91.080 ;
    END
  END core0_data_print[13]
  PIN core0_data_print[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 97.280 400.000 97.880 ;
    END
  END core0_data_print[14]
  PIN core0_data_print[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 101.360 400.000 101.960 ;
    END
  END core0_data_print[15]
  PIN core0_data_print[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END core0_data_print[16]
  PIN core0_data_print[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 114.280 400.000 114.880 ;
    END
  END core0_data_print[17]
  PIN core0_data_print[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END core0_data_print[18]
  PIN core0_data_print[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 130.600 400.000 131.200 ;
    END
  END core0_data_print[19]
  PIN core0_data_print[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 11.600 400.000 12.200 ;
    END
  END core0_data_print[1]
  PIN core0_data_print[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END core0_data_print[20]
  PIN core0_data_print[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 396.000 132.850 400.000 ;
    END
  END core0_data_print[21]
  PIN core0_data_print[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END core0_data_print[22]
  PIN core0_data_print[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END core0_data_print[23]
  PIN core0_data_print[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 146.920 400.000 147.520 ;
    END
  END core0_data_print[24]
  PIN core0_data_print[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 156.440 400.000 157.040 ;
    END
  END core0_data_print[25]
  PIN core0_data_print[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END core0_data_print[26]
  PIN core0_data_print[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 396.000 165.050 400.000 ;
    END
  END core0_data_print[27]
  PIN core0_data_print[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END core0_data_print[28]
  PIN core0_data_print[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END core0_data_print[29]
  PIN core0_data_print[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END core0_data_print[2]
  PIN core0_data_print[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END core0_data_print[30]
  PIN core0_data_print[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 194.520 400.000 195.120 ;
    END
  END core0_data_print[31]
  PIN core0_data_print[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 22.480 400.000 23.080 ;
    END
  END core0_data_print[3]
  PIN core0_data_print[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 396.000 27.970 400.000 ;
    END
  END core0_data_print[4]
  PIN core0_data_print[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 396.000 39.470 400.000 ;
    END
  END core0_data_print[5]
  PIN core0_data_print[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END core0_data_print[6]
  PIN core0_data_print[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 396.000 47.290 400.000 ;
    END
  END core0_data_print[7]
  PIN core0_data_print[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END core0_data_print[8]
  PIN core0_data_print[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END core0_data_print[9]
  PIN csb0_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 2.080 400.000 2.680 ;
    END
  END csb0_to_sram
  PIN data_out_to_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 396.000 2.210 400.000 ;
    END
  END data_out_to_core[0]
  PIN data_out_to_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END data_out_to_core[10]
  PIN data_out_to_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END data_out_to_core[11]
  PIN data_out_to_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 83.000 400.000 83.600 ;
    END
  END data_out_to_core[12]
  PIN data_out_to_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 91.840 400.000 92.440 ;
    END
  END data_out_to_core[13]
  PIN data_out_to_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END data_out_to_core[14]
  PIN data_out_to_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 396.000 94.210 400.000 ;
    END
  END data_out_to_core[15]
  PIN data_out_to_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 396.000 98.810 400.000 ;
    END
  END data_out_to_core[16]
  PIN data_out_to_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 115.640 400.000 116.240 ;
    END
  END data_out_to_core[17]
  PIN data_out_to_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 396.000 108.930 400.000 ;
    END
  END data_out_to_core[18]
  PIN data_out_to_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END data_out_to_core[19]
  PIN data_out_to_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END data_out_to_core[1]
  PIN data_out_to_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 396.000 123.190 400.000 ;
    END
  END data_out_to_core[20]
  PIN data_out_to_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END data_out_to_core[21]
  PIN data_out_to_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 139.440 400.000 140.040 ;
    END
  END data_out_to_core[22]
  PIN data_out_to_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 396.000 144.350 400.000 ;
    END
  END data_out_to_core[23]
  PIN data_out_to_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END data_out_to_core[24]
  PIN data_out_to_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 157.800 400.000 158.400 ;
    END
  END data_out_to_core[25]
  PIN data_out_to_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 161.880 400.000 162.480 ;
    END
  END data_out_to_core[26]
  PIN data_out_to_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END data_out_to_core[27]
  PIN data_out_to_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 174.800 400.000 175.400 ;
    END
  END data_out_to_core[28]
  PIN data_out_to_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 396.000 171.490 400.000 ;
    END
  END data_out_to_core[29]
  PIN data_out_to_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 17.040 400.000 17.640 ;
    END
  END data_out_to_core[2]
  PIN data_out_to_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END data_out_to_core[30]
  PIN data_out_to_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 396.000 179.770 400.000 ;
    END
  END data_out_to_core[31]
  PIN data_out_to_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 24.520 400.000 25.120 ;
    END
  END data_out_to_core[3]
  PIN data_out_to_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 27.920 400.000 28.520 ;
    END
  END data_out_to_core[4]
  PIN data_out_to_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END data_out_to_core[5]
  PIN data_out_to_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END data_out_to_core[6]
  PIN data_out_to_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END data_out_to_core[7]
  PIN data_out_to_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 49.680 400.000 50.280 ;
    END
  END data_out_to_core[8]
  PIN data_out_to_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 59.200 400.000 59.800 ;
    END
  END data_out_to_core[9]
  PIN data_to_core_mem[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 6.160 400.000 6.760 ;
    END
  END data_to_core_mem[0]
  PIN data_to_core_mem[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END data_to_core_mem[10]
  PIN data_to_core_mem[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END data_to_core_mem[11]
  PIN data_to_core_mem[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END data_to_core_mem[12]
  PIN data_to_core_mem[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 93.880 400.000 94.480 ;
    END
  END data_to_core_mem[13]
  PIN data_to_core_mem[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 396.000 89.150 400.000 ;
    END
  END data_to_core_mem[14]
  PIN data_to_core_mem[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END data_to_core_mem[15]
  PIN data_to_core_mem[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END data_to_core_mem[16]
  PIN data_to_core_mem[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 117.680 400.000 118.280 ;
    END
  END data_to_core_mem[17]
  PIN data_to_core_mem[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END data_to_core_mem[18]
  PIN data_to_core_mem[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END data_to_core_mem[19]
  PIN data_to_core_mem[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 396.000 7.270 400.000 ;
    END
  END data_to_core_mem[1]
  PIN data_to_core_mem[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END data_to_core_mem[20]
  PIN data_to_core_mem[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END data_to_core_mem[21]
  PIN data_to_core_mem[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END data_to_core_mem[22]
  PIN data_to_core_mem[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END data_to_core_mem[23]
  PIN data_to_core_mem[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 148.960 400.000 149.560 ;
    END
  END data_to_core_mem[24]
  PIN data_to_core_mem[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 396.000 157.230 400.000 ;
    END
  END data_to_core_mem[25]
  PIN data_to_core_mem[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 163.920 400.000 164.520 ;
    END
  END data_to_core_mem[26]
  PIN data_to_core_mem[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END data_to_core_mem[27]
  PIN data_to_core_mem[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END data_to_core_mem[28]
  PIN data_to_core_mem[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END data_to_core_mem[29]
  PIN data_to_core_mem[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END data_to_core_mem[2]
  PIN data_to_core_mem[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END data_to_core_mem[30]
  PIN data_to_core_mem[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END data_to_core_mem[31]
  PIN data_to_core_mem[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END data_to_core_mem[3]
  PIN data_to_core_mem[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 396.000 29.810 400.000 ;
    END
  END data_to_core_mem[4]
  PIN data_to_core_mem[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END data_to_core_mem[5]
  PIN data_to_core_mem[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END data_to_core_mem[6]
  PIN data_to_core_mem[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END data_to_core_mem[7]
  PIN data_to_core_mem[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 396.000 53.730 400.000 ;
    END
  END data_to_core_mem[8]
  PIN data_to_core_mem[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 61.240 400.000 61.840 ;
    END
  END data_to_core_mem[9]
  PIN din0_to_sram[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END din0_to_sram[0]
  PIN din0_to_sram[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 396.000 66.610 400.000 ;
    END
  END din0_to_sram[10]
  PIN din0_to_sram[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 73.480 400.000 74.080 ;
    END
  END din0_to_sram[11]
  PIN din0_to_sram[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 396.000 76.270 400.000 ;
    END
  END din0_to_sram[12]
  PIN din0_to_sram[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END din0_to_sram[13]
  PIN din0_to_sram[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END din0_to_sram[14]
  PIN din0_to_sram[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END din0_to_sram[15]
  PIN din0_to_sram[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 108.840 400.000 109.440 ;
    END
  END din0_to_sram[16]
  PIN din0_to_sram[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END din0_to_sram[17]
  PIN din0_to_sram[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 121.760 400.000 122.360 ;
    END
  END din0_to_sram[18]
  PIN din0_to_sram[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END din0_to_sram[19]
  PIN din0_to_sram[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END din0_to_sram[1]
  PIN din0_to_sram[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END din0_to_sram[20]
  PIN din0_to_sram[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END din0_to_sram[21]
  PIN din0_to_sram[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END din0_to_sram[22]
  PIN din0_to_sram[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 396.000 145.730 400.000 ;
    END
  END din0_to_sram[23]
  PIN din0_to_sram[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END din0_to_sram[24]
  PIN din0_to_sram[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 396.000 158.610 400.000 ;
    END
  END din0_to_sram[25]
  PIN din0_to_sram[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END din0_to_sram[26]
  PIN din0_to_sram[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 396.000 166.890 400.000 ;
    END
  END din0_to_sram[27]
  PIN din0_to_sram[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 176.160 400.000 176.760 ;
    END
  END din0_to_sram[28]
  PIN din0_to_sram[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END din0_to_sram[29]
  PIN din0_to_sram[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 396.000 18.310 400.000 ;
    END
  END din0_to_sram[2]
  PIN din0_to_sram[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 396.000 174.710 400.000 ;
    END
  END din0_to_sram[30]
  PIN din0_to_sram[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 196.560 400.000 197.160 ;
    END
  END din0_to_sram[31]
  PIN din0_to_sram[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END din0_to_sram[3]
  PIN din0_to_sram[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 396.000 31.190 400.000 ;
    END
  END din0_to_sram[4]
  PIN din0_to_sram[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 33.360 400.000 33.960 ;
    END
  END din0_to_sram[5]
  PIN din0_to_sram[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 40.840 400.000 41.440 ;
    END
  END din0_to_sram[6]
  PIN din0_to_sram[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 396.000 49.130 400.000 ;
    END
  END din0_to_sram[7]
  PIN din0_to_sram[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 51.720 400.000 52.320 ;
    END
  END din0_to_sram[8]
  PIN din0_to_sram[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END din0_to_sram[9]
  PIN dout0_to_sram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END dout0_to_sram[0]
  PIN dout0_to_sram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.040 400.000 68.640 ;
    END
  END dout0_to_sram[10]
  PIN dout0_to_sram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END dout0_to_sram[11]
  PIN dout0_to_sram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END dout0_to_sram[12]
  PIN dout0_to_sram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END dout0_to_sram[13]
  PIN dout0_to_sram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END dout0_to_sram[14]
  PIN dout0_to_sram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 103.400 400.000 104.000 ;
    END
  END dout0_to_sram[15]
  PIN dout0_to_sram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 396.000 100.650 400.000 ;
    END
  END dout0_to_sram[16]
  PIN dout0_to_sram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 396.000 103.870 400.000 ;
    END
  END dout0_to_sram[17]
  PIN dout0_to_sram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 396.000 110.310 400.000 ;
    END
  END dout0_to_sram[18]
  PIN dout0_to_sram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 396.000 116.750 400.000 ;
    END
  END dout0_to_sram[19]
  PIN dout0_to_sram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 396.000 8.650 400.000 ;
    END
  END dout0_to_sram[1]
  PIN dout0_to_sram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END dout0_to_sram[20]
  PIN dout0_to_sram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 396.000 134.690 400.000 ;
    END
  END dout0_to_sram[21]
  PIN dout0_to_sram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 396.000 139.290 400.000 ;
    END
  END dout0_to_sram[22]
  PIN dout0_to_sram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END dout0_to_sram[23]
  PIN dout0_to_sram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 151.000 400.000 151.600 ;
    END
  END dout0_to_sram[24]
  PIN dout0_to_sram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END dout0_to_sram[25]
  PIN dout0_to_sram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END dout0_to_sram[26]
  PIN dout0_to_sram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END dout0_to_sram[27]
  PIN dout0_to_sram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END dout0_to_sram[28]
  PIN dout0_to_sram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 183.640 400.000 184.240 ;
    END
  END dout0_to_sram[29]
  PIN dout0_to_sram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END dout0_to_sram[2]
  PIN dout0_to_sram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 396.000 176.550 400.000 ;
    END
  END dout0_to_sram[30]
  PIN dout0_to_sram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END dout0_to_sram[31]
  PIN dout0_to_sram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END dout0_to_sram[3]
  PIN dout0_to_sram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END dout0_to_sram[4]
  PIN dout0_to_sram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END dout0_to_sram[5]
  PIN dout0_to_sram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END dout0_to_sram[6]
  PIN dout0_to_sram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 44.240 400.000 44.840 ;
    END
  END dout0_to_sram[7]
  PIN dout0_to_sram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 53.760 400.000 54.360 ;
    END
  END dout0_to_sram[8]
  PIN dout0_to_sram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END dout0_to_sram[9]
  PIN is_loading_memory_into_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END is_loading_memory_into_core
  PIN is_ready_dataout_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END is_ready_dataout_core0
  PIN is_ready_print_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END is_ready_print_core0
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 396.000 345.830 400.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 335.960 400.000 336.560 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 396.000 350.890 400.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 356.360 400.000 356.960 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 396.000 358.710 400.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 361.800 400.000 362.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 365.200 400.000 365.800 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 370.640 400.000 371.240 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 396.000 370.210 400.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 396.000 378.030 400.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 396.000 384.470 400.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 396.000 389.530 400.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 396.000 394.130 400.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 398.520 400.000 399.120 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 396.000 78.110 400.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 396.000 84.550 400.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 99.320 400.000 99.920 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 396.000 125.030 400.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 136.040 400.000 136.640 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 396.000 147.570 400.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 152.360 400.000 152.960 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 18.400 400.000 19.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 396.000 177.930 400.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 396.000 182.990 400.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 396.000 187.590 400.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 396.000 195.870 400.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 396.000 199.090 400.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 396.000 202.310 400.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.920 400.000 215.520 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 396.000 207.370 400.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 396.000 215.190 400.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 396.000 229.910 400.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 29.960 400.000 30.560 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 229.880 400.000 230.480 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 396.000 239.570 400.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 396.000 240.950 400.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 242.800 400.000 243.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 396.000 255.670 400.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 396.000 263.490 400.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 396.000 276.370 400.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 266.600 400.000 267.200 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 396.000 40.850 400.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 396.000 289.250 400.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 275.440 400.000 276.040 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.840 400.000 279.440 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 396.000 302.590 400.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 288.360 400.000 288.960 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 396.000 316.850 400.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 301.280 400.000 301.880 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 396.000 321.910 400.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 308.760 400.000 309.360 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 396.000 55.570 400.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 396.000 332.950 400.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 323.040 400.000 323.640 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.920 400.000 334.520 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 396.000 349.050 400.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 343.440 400.000 344.040 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 348.880 400.000 349.480 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 396.000 352.270 400.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 363.840 400.000 364.440 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 396.000 361.930 400.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 372.680 400.000 373.280 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 396.000 365.150 400.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 396.000 371.590 400.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 396.000 374.810 400.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 396.000 376.650 400.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 396.000 379.870 400.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 393.080 400.000 393.680 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 394.440 400.000 395.040 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 396.000 397.350 400.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 396.000 79.490 400.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 396.000 90.990 400.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 396.000 95.590 400.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.120 400.000 123.720 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 396.000 10.490 400.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 396.000 126.410 400.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 396.000 141.130 400.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 396.000 152.170 400.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 20.440 400.000 21.040 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 189.080 400.000 189.680 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 198.600 400.000 199.200 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 396.000 184.370 400.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 202.000 400.000 202.600 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 396.000 197.250 400.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 396.000 204.150 400.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 396.000 205.530 400.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 396.000 208.750 400.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 220.360 400.000 220.960 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 396.000 221.630 400.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 396.000 231.290 400.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 396.000 236.350 400.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.720 400.000 239.320 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 244.160 400.000 244.760 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 396.000 260.270 400.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 35.400 400.000 36.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 249.600 400.000 250.200 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 396.000 265.330 400.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 396.000 274.990 400.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 396.000 278.210 400.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 396.000 282.810 400.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 396.000 42.690 400.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 396.000 287.870 400.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 273.400 400.000 274.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 396.000 292.470 400.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 396.000 298.910 400.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 282.920 400.000 283.520 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 293.800 400.000 294.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 396.000 323.290 400.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 396.000 329.730 400.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 55.120 400.000 55.720 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 396.000 331.570 400.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 312.160 400.000 312.760 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 315.560 400.000 316.160 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 317.600 400.000 318.200 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 327.120 400.000 327.720 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 62.600 400.000 63.200 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 7.520 400.000 8.120 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 396.000 347.670 400.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 339.360 400.000 339.960 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 341.400 400.000 342.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 350.920 400.000 351.520 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 396.000 355.490 400.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.000 4.000 372.600 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 396.000 363.770 400.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 376.080 400.000 376.680 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 380.160 400.000 380.760 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 396.000 69.830 400.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 385.600 400.000 386.200 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 396.000 381.250 400.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 396.000 386.310 400.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 396.000 390.910 400.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 396.000 392.750 400.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 396.480 400.000 397.080 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 104.760 400.000 105.360 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 396.000 102.490 400.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 119.720 400.000 120.320 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 125.160 400.000 125.760 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 396.000 11.870 400.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 396.000 128.250 400.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 138.080 400.000 138.680 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 141.480 400.000 142.080 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 396.000 154.010 400.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.840 400.000 160.440 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 396.000 163.670 400.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 396.000 168.270 400.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 178.200 400.000 178.800 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 396.000 173.330 400.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 396.000 186.210 400.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 396.000 190.810 400.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.040 400.000 204.640 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 0.000 217.030 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 396.000 23.370 400.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 396.000 210.590 400.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.960 400.000 217.560 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 396.000 217.030 400.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 396.000 223.470 400.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 224.440 400.000 225.040 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 396.000 234.510 400.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 396.000 33.030 400.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 233.280 400.000 233.880 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 396.000 242.790 400.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 396.000 247.390 400.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 396.000 250.610 400.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 396.000 269.930 400.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 255.040 400.000 255.640 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 262.520 400.000 263.120 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 396.000 279.590 400.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 270.000 400.000 270.600 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 277.480 400.000 278.080 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 396.000 294.310 400.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 396.000 300.750 400.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 396.000 50.510 400.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 396.000 307.190 400.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 297.200 400.000 297.800 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 299.240 400.000 299.840 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 396.000 320.070 400.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 396.000 325.130 400.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 396.000 326.510 400.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 396.000 56.950 400.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 310.120 400.000 310.720 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 396.000 334.790 400.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 319.640 400.000 320.240 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 325.080 400.000 325.680 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 328.480 400.000 329.080 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 64.640 400.000 65.240 ;
    END
  END la_oenb[9]
  PIN rd_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 396.000 4.050 400.000 ;
    END
  END rd_data_out[0]
  PIN rd_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END rd_data_out[100]
  PIN rd_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 338.000 400.000 338.600 ;
    END
  END rd_data_out[101]
  PIN rd_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END rd_data_out[102]
  PIN rd_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END rd_data_out[103]
  PIN rd_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END rd_data_out[104]
  PIN rd_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END rd_data_out[105]
  PIN rd_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 352.280 400.000 352.880 ;
    END
  END rd_data_out[106]
  PIN rd_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END rd_data_out[107]
  PIN rd_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.720 400.000 358.320 ;
    END
  END rd_data_out[108]
  PIN rd_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 396.000 360.550 400.000 ;
    END
  END rd_data_out[109]
  PIN rd_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END rd_data_out[10]
  PIN rd_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END rd_data_out[110]
  PIN rd_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END rd_data_out[111]
  PIN rd_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END rd_data_out[112]
  PIN rd_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END rd_data_out[113]
  PIN rd_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 367.240 400.000 367.840 ;
    END
  END rd_data_out[114]
  PIN rd_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END rd_data_out[115]
  PIN rd_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 396.000 366.990 400.000 ;
    END
  END rd_data_out[116]
  PIN rd_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 378.120 400.000 378.720 ;
    END
  END rd_data_out[117]
  PIN rd_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 396.000 373.430 400.000 ;
    END
  END rd_data_out[118]
  PIN rd_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END rd_data_out[119]
  PIN rd_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 75.520 400.000 76.120 ;
    END
  END rd_data_out[11]
  PIN rd_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 387.640 400.000 388.240 ;
    END
  END rd_data_out[120]
  PIN rd_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 391.040 400.000 391.640 ;
    END
  END rd_data_out[121]
  PIN rd_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 396.000 387.690 400.000 ;
    END
  END rd_data_out[122]
  PIN rd_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END rd_data_out[123]
  PIN rd_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END rd_data_out[124]
  PIN rd_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END rd_data_out[125]
  PIN rd_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END rd_data_out[126]
  PIN rd_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END rd_data_out[127]
  PIN rd_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 396.000 81.330 400.000 ;
    END
  END rd_data_out[12]
  PIN rd_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END rd_data_out[13]
  PIN rd_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END rd_data_out[14]
  PIN rd_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END rd_data_out[15]
  PIN rd_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END rd_data_out[16]
  PIN rd_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END rd_data_out[17]
  PIN rd_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END rd_data_out[18]
  PIN rd_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 396.000 118.590 400.000 ;
    END
  END rd_data_out[19]
  PIN rd_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 396.000 13.710 400.000 ;
    END
  END rd_data_out[1]
  PIN rd_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END rd_data_out[20]
  PIN rd_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END rd_data_out[21]
  PIN rd_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 396.000 142.510 400.000 ;
    END
  END rd_data_out[22]
  PIN rd_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 143.520 400.000 144.120 ;
    END
  END rd_data_out[23]
  PIN rd_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 154.400 400.000 155.000 ;
    END
  END rd_data_out[24]
  PIN rd_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END rd_data_out[25]
  PIN rd_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 165.280 400.000 165.880 ;
    END
  END rd_data_out[26]
  PIN rd_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.720 400.000 171.320 ;
    END
  END rd_data_out[27]
  PIN rd_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END rd_data_out[28]
  PIN rd_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 185.680 400.000 186.280 ;
    END
  END rd_data_out[29]
  PIN rd_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END rd_data_out[2]
  PIN rd_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END rd_data_out[30]
  PIN rd_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END rd_data_out[31]
  PIN rd_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END rd_data_out[32]
  PIN rd_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END rd_data_out[33]
  PIN rd_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 396.000 192.650 400.000 ;
    END
  END rd_data_out[34]
  PIN rd_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END rd_data_out[35]
  PIN rd_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 206.080 400.000 206.680 ;
    END
  END rd_data_out[36]
  PIN rd_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 396.000 200.930 400.000 ;
    END
  END rd_data_out[37]
  PIN rd_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 211.520 400.000 212.120 ;
    END
  END rd_data_out[38]
  PIN rd_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 212.880 400.000 213.480 ;
    END
  END rd_data_out[39]
  PIN rd_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 396.000 24.750 400.000 ;
    END
  END rd_data_out[3]
  PIN rd_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END rd_data_out[40]
  PIN rd_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END rd_data_out[41]
  PIN rd_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 396.000 211.970 400.000 ;
    END
  END rd_data_out[42]
  PIN rd_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 396.000 213.810 400.000 ;
    END
  END rd_data_out[43]
  PIN rd_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 396.000 218.410 400.000 ;
    END
  END rd_data_out[44]
  PIN rd_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 222.400 400.000 223.000 ;
    END
  END rd_data_out[45]
  PIN rd_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 396.000 224.850 400.000 ;
    END
  END rd_data_out[46]
  PIN rd_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 396.000 226.690 400.000 ;
    END
  END rd_data_out[47]
  PIN rd_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 225.800 400.000 226.400 ;
    END
  END rd_data_out[48]
  PIN rd_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.840 400.000 228.440 ;
    END
  END rd_data_out[49]
  PIN rd_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END rd_data_out[4]
  PIN rd_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 396.000 237.730 400.000 ;
    END
  END rd_data_out[50]
  PIN rd_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END rd_data_out[51]
  PIN rd_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END rd_data_out[52]
  PIN rd_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END rd_data_out[53]
  PIN rd_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 240.760 400.000 241.360 ;
    END
  END rd_data_out[54]
  PIN rd_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 396.000 249.230 400.000 ;
    END
  END rd_data_out[55]
  PIN rd_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 396.000 252.450 400.000 ;
    END
  END rd_data_out[56]
  PIN rd_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 246.200 400.000 246.800 ;
    END
  END rd_data_out[57]
  PIN rd_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 396.000 257.050 400.000 ;
    END
  END rd_data_out[58]
  PIN rd_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 396.000 262.110 400.000 ;
    END
  END rd_data_out[59]
  PIN rd_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END rd_data_out[5]
  PIN rd_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END rd_data_out[60]
  PIN rd_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 396.000 266.710 400.000 ;
    END
  END rd_data_out[61]
  PIN rd_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 251.640 400.000 252.240 ;
    END
  END rd_data_out[62]
  PIN rd_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 257.080 400.000 257.680 ;
    END
  END rd_data_out[63]
  PIN rd_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 259.120 400.000 259.720 ;
    END
  END rd_data_out[64]
  PIN rd_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 261.160 400.000 261.760 ;
    END
  END rd_data_out[65]
  PIN rd_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END rd_data_out[66]
  PIN rd_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 396.000 281.430 400.000 ;
    END
  END rd_data_out[67]
  PIN rd_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END rd_data_out[68]
  PIN rd_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 396.000 284.650 400.000 ;
    END
  END rd_data_out[69]
  PIN rd_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END rd_data_out[6]
  PIN rd_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END rd_data_out[70]
  PIN rd_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 272.040 400.000 272.640 ;
    END
  END rd_data_out[71]
  PIN rd_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END rd_data_out[72]
  PIN rd_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END rd_data_out[73]
  PIN rd_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 396.000 295.690 400.000 ;
    END
  END rd_data_out[74]
  PIN rd_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 396.000 297.530 400.000 ;
    END
  END rd_data_out[75]
  PIN rd_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 280.880 400.000 281.480 ;
    END
  END rd_data_out[76]
  PIN rd_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 396.000 303.970 400.000 ;
    END
  END rd_data_out[77]
  PIN rd_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 286.320 400.000 286.920 ;
    END
  END rd_data_out[78]
  PIN rd_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 290.400 400.000 291.000 ;
    END
  END rd_data_out[79]
  PIN rd_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 396.000 52.350 400.000 ;
    END
  END rd_data_out[7]
  PIN rd_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 396.000 309.030 400.000 ;
    END
  END rd_data_out[80]
  PIN rd_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 295.840 400.000 296.440 ;
    END
  END rd_data_out[81]
  PIN rd_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 396.000 313.630 400.000 ;
    END
  END rd_data_out[82]
  PIN rd_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 396.000 318.690 400.000 ;
    END
  END rd_data_out[83]
  PIN rd_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END rd_data_out[84]
  PIN rd_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END rd_data_out[85]
  PIN rd_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END rd_data_out[86]
  PIN rd_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 303.320 400.000 303.920 ;
    END
  END rd_data_out[87]
  PIN rd_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.720 400.000 307.320 ;
    END
  END rd_data_out[88]
  PIN rd_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END rd_data_out[89]
  PIN rd_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END rd_data_out[8]
  PIN rd_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END rd_data_out[90]
  PIN rd_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 314.200 400.000 314.800 ;
    END
  END rd_data_out[91]
  PIN rd_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 396.000 336.170 400.000 ;
    END
  END rd_data_out[92]
  PIN rd_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 396.000 338.010 400.000 ;
    END
  END rd_data_out[93]
  PIN rd_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.680 400.000 322.280 ;
    END
  END rd_data_out[94]
  PIN rd_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 396.000 341.230 400.000 ;
    END
  END rd_data_out[95]
  PIN rd_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END rd_data_out[96]
  PIN rd_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END rd_data_out[97]
  PIN rd_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 330.520 400.000 331.120 ;
    END
  END rd_data_out[98]
  PIN rd_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 332.560 400.000 333.160 ;
    END
  END rd_data_out[99]
  PIN rd_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 66.680 400.000 67.280 ;
    END
  END rd_data_out[9]
  PIN read_enable_to_Elpis
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END read_enable_to_Elpis
  PIN read_interactive_req_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END read_interactive_req_core0
  PIN read_value_to_Elpis[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END read_value_to_Elpis[0]
  PIN read_value_to_Elpis[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END read_value_to_Elpis[10]
  PIN read_value_to_Elpis[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 77.560 400.000 78.160 ;
    END
  END read_value_to_Elpis[11]
  PIN read_value_to_Elpis[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 396.000 82.710 400.000 ;
    END
  END read_value_to_Elpis[12]
  PIN read_value_to_Elpis[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 396.000 85.930 400.000 ;
    END
  END read_value_to_Elpis[13]
  PIN read_value_to_Elpis[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END read_value_to_Elpis[14]
  PIN read_value_to_Elpis[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 106.800 400.000 107.400 ;
    END
  END read_value_to_Elpis[15]
  PIN read_value_to_Elpis[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 110.200 400.000 110.800 ;
    END
  END read_value_to_Elpis[16]
  PIN read_value_to_Elpis[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END read_value_to_Elpis[17]
  PIN read_value_to_Elpis[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 396.000 112.150 400.000 ;
    END
  END read_value_to_Elpis[18]
  PIN read_value_to_Elpis[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 132.640 400.000 133.240 ;
    END
  END read_value_to_Elpis[19]
  PIN read_value_to_Elpis[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 396.000 15.090 400.000 ;
    END
  END read_value_to_Elpis[1]
  PIN read_value_to_Elpis[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 134.000 400.000 134.600 ;
    END
  END read_value_to_Elpis[20]
  PIN read_value_to_Elpis[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END read_value_to_Elpis[21]
  PIN read_value_to_Elpis[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END read_value_to_Elpis[22]
  PIN read_value_to_Elpis[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 396.000 148.950 400.000 ;
    END
  END read_value_to_Elpis[23]
  PIN read_value_to_Elpis[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 396.000 155.390 400.000 ;
    END
  END read_value_to_Elpis[24]
  PIN read_value_to_Elpis[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 396.000 160.450 400.000 ;
    END
  END read_value_to_Elpis[25]
  PIN read_value_to_Elpis[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END read_value_to_Elpis[26]
  PIN read_value_to_Elpis[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 172.760 400.000 173.360 ;
    END
  END read_value_to_Elpis[27]
  PIN read_value_to_Elpis[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.240 400.000 180.840 ;
    END
  END read_value_to_Elpis[28]
  PIN read_value_to_Elpis[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 187.720 400.000 188.320 ;
    END
  END read_value_to_Elpis[29]
  PIN read_value_to_Elpis[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END read_value_to_Elpis[2]
  PIN read_value_to_Elpis[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 191.120 400.000 191.720 ;
    END
  END read_value_to_Elpis[30]
  PIN read_value_to_Elpis[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 200.640 400.000 201.240 ;
    END
  END read_value_to_Elpis[31]
  PIN read_value_to_Elpis[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END read_value_to_Elpis[3]
  PIN read_value_to_Elpis[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 31.320 400.000 31.920 ;
    END
  END read_value_to_Elpis[4]
  PIN read_value_to_Elpis[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END read_value_to_Elpis[5]
  PIN read_value_to_Elpis[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 396.000 44.070 400.000 ;
    END
  END read_value_to_Elpis[6]
  PIN read_value_to_Elpis[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END read_value_to_Elpis[7]
  PIN read_value_to_Elpis[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 396.000 58.790 400.000 ;
    END
  END read_value_to_Elpis[8]
  PIN read_value_to_Elpis[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END read_value_to_Elpis[9]
  PIN ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END ready
  PIN req_out_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END req_out_core0
  PIN requested
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END requested
  PIN reset_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END reset_core
  PIN reset_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END reset_mem_req
  PIN rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END rst
  PIN spare_wen0_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 4.120 400.000 4.720 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_rst_i
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 396.000 68.450 400.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 85.040 400.000 85.640 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.920 400.000 96.520 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 396.000 105.710 400.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 127.200 400.000 127.800 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 396.000 119.970 400.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 12.960 400.000 13.560 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 396.000 129.630 400.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 396.000 136.070 400.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 396.000 150.790 400.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 167.320 400.000 167.920 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 182.280 400.000 182.880 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 396.000 20.150 400.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 396.000 34.410 400.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 396.000 60.170 400.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END wbs_dat_o[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END we
  PIN we_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 0.720 400.000 1.320 ;
    END
  END we_to_sram
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 396.000 5.430 400.000 ;
    END
  END wr_data[0]
  PIN wr_data[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END wr_data[100]
  PIN wr_data[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END wr_data[101]
  PIN wr_data[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.520 4.000 348.120 ;
    END
  END wr_data[102]
  PIN wr_data[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END wr_data[103]
  PIN wr_data[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 345.480 400.000 346.080 ;
    END
  END wr_data[104]
  PIN wr_data[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 346.840 400.000 347.440 ;
    END
  END wr_data[105]
  PIN wr_data[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 354.320 400.000 354.920 ;
    END
  END wr_data[106]
  PIN wr_data[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 396.000 354.110 400.000 ;
    END
  END wr_data[107]
  PIN wr_data[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 396.000 357.330 400.000 ;
    END
  END wr_data[108]
  PIN wr_data[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END wr_data[109]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 70.080 400.000 70.680 ;
    END
  END wr_data[10]
  PIN wr_data[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 359.760 400.000 360.360 ;
    END
  END wr_data[110]
  PIN wr_data[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END wr_data[111]
  PIN wr_data[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END wr_data[112]
  PIN wr_data[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END wr_data[113]
  PIN wr_data[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 369.280 400.000 369.880 ;
    END
  END wr_data[114]
  PIN wr_data[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 374.720 400.000 375.320 ;
    END
  END wr_data[115]
  PIN wr_data[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 396.000 368.370 400.000 ;
    END
  END wr_data[116]
  PIN wr_data[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END wr_data[117]
  PIN wr_data[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 382.200 400.000 382.800 ;
    END
  END wr_data[118]
  PIN wr_data[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 383.560 400.000 384.160 ;
    END
  END wr_data[119]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 78.920 400.000 79.520 ;
    END
  END wr_data[11]
  PIN wr_data[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 389.000 400.000 389.600 ;
    END
  END wr_data[120]
  PIN wr_data[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 396.000 383.090 400.000 ;
    END
  END wr_data[121]
  PIN wr_data[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END wr_data[122]
  PIN wr_data[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END wr_data[123]
  PIN wr_data[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END wr_data[124]
  PIN wr_data[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 396.000 395.970 400.000 ;
    END
  END wr_data[125]
  PIN wr_data[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 396.000 399.190 400.000 ;
    END
  END wr_data[126]
  PIN wr_data[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END wr_data[127]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wr_data[12]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END wr_data[13]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END wr_data[14]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 396.000 97.430 400.000 ;
    END
  END wr_data[15]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.240 400.000 112.840 ;
    END
  END wr_data[16]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wr_data[17]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 396.000 113.530 400.000 ;
    END
  END wr_data[18]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 396.000 121.810 400.000 ;
    END
  END wr_data[19]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END wr_data[1]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 396.000 131.470 400.000 ;
    END
  END wr_data[20]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 396.000 137.910 400.000 ;
    END
  END wr_data[21]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wr_data[22]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 145.560 400.000 146.160 ;
    END
  END wr_data[23]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wr_data[24]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 396.000 161.830 400.000 ;
    END
  END wr_data[25]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 169.360 400.000 169.960 ;
    END
  END wr_data[26]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 396.000 170.110 400.000 ;
    END
  END wr_data[27]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END wr_data[28]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END wr_data[29]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 396.000 21.530 400.000 ;
    END
  END wr_data[2]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.160 400.000 193.760 ;
    END
  END wr_data[30]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 396.000 181.150 400.000 ;
    END
  END wr_data[31]
  PIN wr_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END wr_data[32]
  PIN wr_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 396.000 189.430 400.000 ;
    END
  END wr_data[33]
  PIN wr_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 396.000 194.030 400.000 ;
    END
  END wr_data[34]
  PIN wr_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wr_data[35]
  PIN wr_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 207.440 400.000 208.040 ;
    END
  END wr_data[36]
  PIN wr_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 209.480 400.000 210.080 ;
    END
  END wr_data[37]
  PIN wr_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END wr_data[38]
  PIN wr_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END wr_data[39]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wr_data[3]
  PIN wr_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END wr_data[40]
  PIN wr_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END wr_data[41]
  PIN wr_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END wr_data[42]
  PIN wr_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END wr_data[43]
  PIN wr_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 218.320 400.000 218.920 ;
    END
  END wr_data[44]
  PIN wr_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 396.000 220.250 400.000 ;
    END
  END wr_data[45]
  PIN wr_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END wr_data[46]
  PIN wr_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 396.000 228.070 400.000 ;
    END
  END wr_data[47]
  PIN wr_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 396.000 233.130 400.000 ;
    END
  END wr_data[48]
  PIN wr_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END wr_data[49]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 396.000 36.250 400.000 ;
    END
  END wr_data[4]
  PIN wr_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 231.240 400.000 231.840 ;
    END
  END wr_data[50]
  PIN wr_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 235.320 400.000 235.920 ;
    END
  END wr_data[51]
  PIN wr_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 236.680 400.000 237.280 ;
    END
  END wr_data[52]
  PIN wr_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 396.000 244.170 400.000 ;
    END
  END wr_data[53]
  PIN wr_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 396.000 246.010 400.000 ;
    END
  END wr_data[54]
  PIN wr_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END wr_data[55]
  PIN wr_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 396.000 253.830 400.000 ;
    END
  END wr_data[56]
  PIN wr_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.240 400.000 248.840 ;
    END
  END wr_data[57]
  PIN wr_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 396.000 258.890 400.000 ;
    END
  END wr_data[58]
  PIN wr_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END wr_data[59]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END wr_data[5]
  PIN wr_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END wr_data[60]
  PIN wr_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 396.000 268.550 400.000 ;
    END
  END wr_data[61]
  PIN wr_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 253.680 400.000 254.280 ;
    END
  END wr_data[62]
  PIN wr_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END wr_data[63]
  PIN wr_data[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 396.000 271.770 400.000 ;
    END
  END wr_data[64]
  PIN wr_data[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 396.000 273.150 400.000 ;
    END
  END wr_data[65]
  PIN wr_data[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 264.560 400.000 265.160 ;
    END
  END wr_data[66]
  PIN wr_data[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END wr_data[67]
  PIN wr_data[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END wr_data[68]
  PIN wr_data[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 267.960 400.000 268.560 ;
    END
  END wr_data[69]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 396.000 45.910 400.000 ;
    END
  END wr_data[6]
  PIN wr_data[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 396.000 286.030 400.000 ;
    END
  END wr_data[70]
  PIN wr_data[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END wr_data[71]
  PIN wr_data[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 396.000 291.090 400.000 ;
    END
  END wr_data[72]
  PIN wr_data[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END wr_data[73]
  PIN wr_data[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END wr_data[74]
  PIN wr_data[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wr_data[75]
  PIN wr_data[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END wr_data[76]
  PIN wr_data[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 284.960 400.000 285.560 ;
    END
  END wr_data[77]
  PIN wr_data[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 396.000 305.810 400.000 ;
    END
  END wr_data[78]
  PIN wr_data[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 291.760 400.000 292.360 ;
    END
  END wr_data[79]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wr_data[7]
  PIN wr_data[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 396.000 310.410 400.000 ;
    END
  END wr_data[80]
  PIN wr_data[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 396.000 312.250 400.000 ;
    END
  END wr_data[81]
  PIN wr_data[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 396.000 315.470 400.000 ;
    END
  END wr_data[82]
  PIN wr_data[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END wr_data[83]
  PIN wr_data[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END wr_data[84]
  PIN wr_data[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END wr_data[85]
  PIN wr_data[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END wr_data[86]
  PIN wr_data[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 304.680 400.000 305.280 ;
    END
  END wr_data[87]
  PIN wr_data[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 396.000 328.350 400.000 ;
    END
  END wr_data[88]
  PIN wr_data[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wr_data[89]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 396.000 62.010 400.000 ;
    END
  END wr_data[8]
  PIN wr_data[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wr_data[90]
  PIN wr_data[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END wr_data[91]
  PIN wr_data[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END wr_data[92]
  PIN wr_data[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END wr_data[93]
  PIN wr_data[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 396.000 339.390 400.000 ;
    END
  END wr_data[94]
  PIN wr_data[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 396.000 342.610 400.000 ;
    END
  END wr_data[95]
  PIN wr_data[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END wr_data[96]
  PIN wr_data[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END wr_data[97]
  PIN wr_data[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END wr_data[98]
  PIN wr_data[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 396.000 344.450 400.000 ;
    END
  END wr_data[99]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wr_data[9]
  OBS
      LAYER li1 ;
        RECT 4.745 10.795 396.835 391.255 ;
      LAYER met1 ;
        RECT 0.530 5.820 399.210 391.300 ;
      LAYER met2 ;
        RECT 1.110 395.720 1.650 399.005 ;
        RECT 2.490 395.720 3.490 399.005 ;
        RECT 4.330 395.720 4.870 399.005 ;
        RECT 5.710 395.720 6.710 399.005 ;
        RECT 7.550 395.720 8.090 399.005 ;
        RECT 8.930 395.720 9.930 399.005 ;
        RECT 10.770 395.720 11.310 399.005 ;
        RECT 12.150 395.720 13.150 399.005 ;
        RECT 13.990 395.720 14.530 399.005 ;
        RECT 15.370 395.720 16.370 399.005 ;
        RECT 17.210 395.720 17.750 399.005 ;
        RECT 18.590 395.720 19.590 399.005 ;
        RECT 20.430 395.720 20.970 399.005 ;
        RECT 21.810 395.720 22.810 399.005 ;
        RECT 23.650 395.720 24.190 399.005 ;
        RECT 25.030 395.720 26.030 399.005 ;
        RECT 26.870 395.720 27.410 399.005 ;
        RECT 28.250 395.720 29.250 399.005 ;
        RECT 30.090 395.720 30.630 399.005 ;
        RECT 31.470 395.720 32.470 399.005 ;
        RECT 33.310 395.720 33.850 399.005 ;
        RECT 34.690 395.720 35.690 399.005 ;
        RECT 36.530 395.720 37.070 399.005 ;
        RECT 37.910 395.720 38.910 399.005 ;
        RECT 39.750 395.720 40.290 399.005 ;
        RECT 41.130 395.720 42.130 399.005 ;
        RECT 42.970 395.720 43.510 399.005 ;
        RECT 44.350 395.720 45.350 399.005 ;
        RECT 46.190 395.720 46.730 399.005 ;
        RECT 47.570 395.720 48.570 399.005 ;
        RECT 49.410 395.720 49.950 399.005 ;
        RECT 50.790 395.720 51.790 399.005 ;
        RECT 52.630 395.720 53.170 399.005 ;
        RECT 54.010 395.720 55.010 399.005 ;
        RECT 55.850 395.720 56.390 399.005 ;
        RECT 57.230 395.720 58.230 399.005 ;
        RECT 59.070 395.720 59.610 399.005 ;
        RECT 60.450 395.720 61.450 399.005 ;
        RECT 62.290 395.720 62.830 399.005 ;
        RECT 63.670 395.720 64.670 399.005 ;
        RECT 65.510 395.720 66.050 399.005 ;
        RECT 66.890 395.720 67.890 399.005 ;
        RECT 68.730 395.720 69.270 399.005 ;
        RECT 70.110 395.720 71.110 399.005 ;
        RECT 71.950 395.720 72.490 399.005 ;
        RECT 73.330 395.720 74.330 399.005 ;
        RECT 75.170 395.720 75.710 399.005 ;
        RECT 76.550 395.720 77.550 399.005 ;
        RECT 78.390 395.720 78.930 399.005 ;
        RECT 79.770 395.720 80.770 399.005 ;
        RECT 81.610 395.720 82.150 399.005 ;
        RECT 82.990 395.720 83.990 399.005 ;
        RECT 84.830 395.720 85.370 399.005 ;
        RECT 86.210 395.720 87.210 399.005 ;
        RECT 88.050 395.720 88.590 399.005 ;
        RECT 89.430 395.720 90.430 399.005 ;
        RECT 91.270 395.720 91.810 399.005 ;
        RECT 92.650 395.720 93.650 399.005 ;
        RECT 94.490 395.720 95.030 399.005 ;
        RECT 95.870 395.720 96.870 399.005 ;
        RECT 97.710 395.720 98.250 399.005 ;
        RECT 99.090 395.720 100.090 399.005 ;
        RECT 100.930 395.720 101.930 399.005 ;
        RECT 102.770 395.720 103.310 399.005 ;
        RECT 104.150 395.720 105.150 399.005 ;
        RECT 105.990 395.720 106.530 399.005 ;
        RECT 107.370 395.720 108.370 399.005 ;
        RECT 109.210 395.720 109.750 399.005 ;
        RECT 110.590 395.720 111.590 399.005 ;
        RECT 112.430 395.720 112.970 399.005 ;
        RECT 113.810 395.720 114.810 399.005 ;
        RECT 115.650 395.720 116.190 399.005 ;
        RECT 117.030 395.720 118.030 399.005 ;
        RECT 118.870 395.720 119.410 399.005 ;
        RECT 120.250 395.720 121.250 399.005 ;
        RECT 122.090 395.720 122.630 399.005 ;
        RECT 123.470 395.720 124.470 399.005 ;
        RECT 125.310 395.720 125.850 399.005 ;
        RECT 126.690 395.720 127.690 399.005 ;
        RECT 128.530 395.720 129.070 399.005 ;
        RECT 129.910 395.720 130.910 399.005 ;
        RECT 131.750 395.720 132.290 399.005 ;
        RECT 133.130 395.720 134.130 399.005 ;
        RECT 134.970 395.720 135.510 399.005 ;
        RECT 136.350 395.720 137.350 399.005 ;
        RECT 138.190 395.720 138.730 399.005 ;
        RECT 139.570 395.720 140.570 399.005 ;
        RECT 141.410 395.720 141.950 399.005 ;
        RECT 142.790 395.720 143.790 399.005 ;
        RECT 144.630 395.720 145.170 399.005 ;
        RECT 146.010 395.720 147.010 399.005 ;
        RECT 147.850 395.720 148.390 399.005 ;
        RECT 149.230 395.720 150.230 399.005 ;
        RECT 151.070 395.720 151.610 399.005 ;
        RECT 152.450 395.720 153.450 399.005 ;
        RECT 154.290 395.720 154.830 399.005 ;
        RECT 155.670 395.720 156.670 399.005 ;
        RECT 157.510 395.720 158.050 399.005 ;
        RECT 158.890 395.720 159.890 399.005 ;
        RECT 160.730 395.720 161.270 399.005 ;
        RECT 162.110 395.720 163.110 399.005 ;
        RECT 163.950 395.720 164.490 399.005 ;
        RECT 165.330 395.720 166.330 399.005 ;
        RECT 167.170 395.720 167.710 399.005 ;
        RECT 168.550 395.720 169.550 399.005 ;
        RECT 170.390 395.720 170.930 399.005 ;
        RECT 171.770 395.720 172.770 399.005 ;
        RECT 173.610 395.720 174.150 399.005 ;
        RECT 174.990 395.720 175.990 399.005 ;
        RECT 176.830 395.720 177.370 399.005 ;
        RECT 178.210 395.720 179.210 399.005 ;
        RECT 180.050 395.720 180.590 399.005 ;
        RECT 181.430 395.720 182.430 399.005 ;
        RECT 183.270 395.720 183.810 399.005 ;
        RECT 184.650 395.720 185.650 399.005 ;
        RECT 186.490 395.720 187.030 399.005 ;
        RECT 187.870 395.720 188.870 399.005 ;
        RECT 189.710 395.720 190.250 399.005 ;
        RECT 191.090 395.720 192.090 399.005 ;
        RECT 192.930 395.720 193.470 399.005 ;
        RECT 194.310 395.720 195.310 399.005 ;
        RECT 196.150 395.720 196.690 399.005 ;
        RECT 197.530 395.720 198.530 399.005 ;
        RECT 199.370 395.720 200.370 399.005 ;
        RECT 201.210 395.720 201.750 399.005 ;
        RECT 202.590 395.720 203.590 399.005 ;
        RECT 204.430 395.720 204.970 399.005 ;
        RECT 205.810 395.720 206.810 399.005 ;
        RECT 207.650 395.720 208.190 399.005 ;
        RECT 209.030 395.720 210.030 399.005 ;
        RECT 210.870 395.720 211.410 399.005 ;
        RECT 212.250 395.720 213.250 399.005 ;
        RECT 214.090 395.720 214.630 399.005 ;
        RECT 215.470 395.720 216.470 399.005 ;
        RECT 217.310 395.720 217.850 399.005 ;
        RECT 218.690 395.720 219.690 399.005 ;
        RECT 220.530 395.720 221.070 399.005 ;
        RECT 221.910 395.720 222.910 399.005 ;
        RECT 223.750 395.720 224.290 399.005 ;
        RECT 225.130 395.720 226.130 399.005 ;
        RECT 226.970 395.720 227.510 399.005 ;
        RECT 228.350 395.720 229.350 399.005 ;
        RECT 230.190 395.720 230.730 399.005 ;
        RECT 231.570 395.720 232.570 399.005 ;
        RECT 233.410 395.720 233.950 399.005 ;
        RECT 234.790 395.720 235.790 399.005 ;
        RECT 236.630 395.720 237.170 399.005 ;
        RECT 238.010 395.720 239.010 399.005 ;
        RECT 239.850 395.720 240.390 399.005 ;
        RECT 241.230 395.720 242.230 399.005 ;
        RECT 243.070 395.720 243.610 399.005 ;
        RECT 244.450 395.720 245.450 399.005 ;
        RECT 246.290 395.720 246.830 399.005 ;
        RECT 247.670 395.720 248.670 399.005 ;
        RECT 249.510 395.720 250.050 399.005 ;
        RECT 250.890 395.720 251.890 399.005 ;
        RECT 252.730 395.720 253.270 399.005 ;
        RECT 254.110 395.720 255.110 399.005 ;
        RECT 255.950 395.720 256.490 399.005 ;
        RECT 257.330 395.720 258.330 399.005 ;
        RECT 259.170 395.720 259.710 399.005 ;
        RECT 260.550 395.720 261.550 399.005 ;
        RECT 262.390 395.720 262.930 399.005 ;
        RECT 263.770 395.720 264.770 399.005 ;
        RECT 265.610 395.720 266.150 399.005 ;
        RECT 266.990 395.720 267.990 399.005 ;
        RECT 268.830 395.720 269.370 399.005 ;
        RECT 270.210 395.720 271.210 399.005 ;
        RECT 272.050 395.720 272.590 399.005 ;
        RECT 273.430 395.720 274.430 399.005 ;
        RECT 275.270 395.720 275.810 399.005 ;
        RECT 276.650 395.720 277.650 399.005 ;
        RECT 278.490 395.720 279.030 399.005 ;
        RECT 279.870 395.720 280.870 399.005 ;
        RECT 281.710 395.720 282.250 399.005 ;
        RECT 283.090 395.720 284.090 399.005 ;
        RECT 284.930 395.720 285.470 399.005 ;
        RECT 286.310 395.720 287.310 399.005 ;
        RECT 288.150 395.720 288.690 399.005 ;
        RECT 289.530 395.720 290.530 399.005 ;
        RECT 291.370 395.720 291.910 399.005 ;
        RECT 292.750 395.720 293.750 399.005 ;
        RECT 294.590 395.720 295.130 399.005 ;
        RECT 295.970 395.720 296.970 399.005 ;
        RECT 297.810 395.720 298.350 399.005 ;
        RECT 299.190 395.720 300.190 399.005 ;
        RECT 301.030 395.720 302.030 399.005 ;
        RECT 302.870 395.720 303.410 399.005 ;
        RECT 304.250 395.720 305.250 399.005 ;
        RECT 306.090 395.720 306.630 399.005 ;
        RECT 307.470 395.720 308.470 399.005 ;
        RECT 309.310 395.720 309.850 399.005 ;
        RECT 310.690 395.720 311.690 399.005 ;
        RECT 312.530 395.720 313.070 399.005 ;
        RECT 313.910 395.720 314.910 399.005 ;
        RECT 315.750 395.720 316.290 399.005 ;
        RECT 317.130 395.720 318.130 399.005 ;
        RECT 318.970 395.720 319.510 399.005 ;
        RECT 320.350 395.720 321.350 399.005 ;
        RECT 322.190 395.720 322.730 399.005 ;
        RECT 323.570 395.720 324.570 399.005 ;
        RECT 325.410 395.720 325.950 399.005 ;
        RECT 326.790 395.720 327.790 399.005 ;
        RECT 328.630 395.720 329.170 399.005 ;
        RECT 330.010 395.720 331.010 399.005 ;
        RECT 331.850 395.720 332.390 399.005 ;
        RECT 333.230 395.720 334.230 399.005 ;
        RECT 335.070 395.720 335.610 399.005 ;
        RECT 336.450 395.720 337.450 399.005 ;
        RECT 338.290 395.720 338.830 399.005 ;
        RECT 339.670 395.720 340.670 399.005 ;
        RECT 341.510 395.720 342.050 399.005 ;
        RECT 342.890 395.720 343.890 399.005 ;
        RECT 344.730 395.720 345.270 399.005 ;
        RECT 346.110 395.720 347.110 399.005 ;
        RECT 347.950 395.720 348.490 399.005 ;
        RECT 349.330 395.720 350.330 399.005 ;
        RECT 351.170 395.720 351.710 399.005 ;
        RECT 352.550 395.720 353.550 399.005 ;
        RECT 354.390 395.720 354.930 399.005 ;
        RECT 355.770 395.720 356.770 399.005 ;
        RECT 357.610 395.720 358.150 399.005 ;
        RECT 358.990 395.720 359.990 399.005 ;
        RECT 360.830 395.720 361.370 399.005 ;
        RECT 362.210 395.720 363.210 399.005 ;
        RECT 364.050 395.720 364.590 399.005 ;
        RECT 365.430 395.720 366.430 399.005 ;
        RECT 367.270 395.720 367.810 399.005 ;
        RECT 368.650 395.720 369.650 399.005 ;
        RECT 370.490 395.720 371.030 399.005 ;
        RECT 371.870 395.720 372.870 399.005 ;
        RECT 373.710 395.720 374.250 399.005 ;
        RECT 375.090 395.720 376.090 399.005 ;
        RECT 376.930 395.720 377.470 399.005 ;
        RECT 378.310 395.720 379.310 399.005 ;
        RECT 380.150 395.720 380.690 399.005 ;
        RECT 381.530 395.720 382.530 399.005 ;
        RECT 383.370 395.720 383.910 399.005 ;
        RECT 384.750 395.720 385.750 399.005 ;
        RECT 386.590 395.720 387.130 399.005 ;
        RECT 387.970 395.720 388.970 399.005 ;
        RECT 389.810 395.720 390.350 399.005 ;
        RECT 391.190 395.720 392.190 399.005 ;
        RECT 393.030 395.720 393.570 399.005 ;
        RECT 394.410 395.720 395.410 399.005 ;
        RECT 396.250 395.720 396.790 399.005 ;
        RECT 397.630 395.720 398.630 399.005 ;
        RECT 0.560 4.280 399.180 395.720 ;
        RECT 1.110 0.835 1.650 4.280 ;
        RECT 2.490 0.835 3.490 4.280 ;
        RECT 4.330 0.835 4.870 4.280 ;
        RECT 5.710 0.835 6.710 4.280 ;
        RECT 7.550 0.835 8.090 4.280 ;
        RECT 8.930 0.835 9.930 4.280 ;
        RECT 10.770 0.835 11.310 4.280 ;
        RECT 12.150 0.835 13.150 4.280 ;
        RECT 13.990 0.835 14.530 4.280 ;
        RECT 15.370 0.835 16.370 4.280 ;
        RECT 17.210 0.835 17.750 4.280 ;
        RECT 18.590 0.835 19.590 4.280 ;
        RECT 20.430 0.835 20.970 4.280 ;
        RECT 21.810 0.835 22.810 4.280 ;
        RECT 23.650 0.835 24.190 4.280 ;
        RECT 25.030 0.835 26.030 4.280 ;
        RECT 26.870 0.835 27.410 4.280 ;
        RECT 28.250 0.835 29.250 4.280 ;
        RECT 30.090 0.835 30.630 4.280 ;
        RECT 31.470 0.835 32.470 4.280 ;
        RECT 33.310 0.835 33.850 4.280 ;
        RECT 34.690 0.835 35.690 4.280 ;
        RECT 36.530 0.835 37.070 4.280 ;
        RECT 37.910 0.835 38.910 4.280 ;
        RECT 39.750 0.835 40.290 4.280 ;
        RECT 41.130 0.835 42.130 4.280 ;
        RECT 42.970 0.835 43.510 4.280 ;
        RECT 44.350 0.835 45.350 4.280 ;
        RECT 46.190 0.835 46.730 4.280 ;
        RECT 47.570 0.835 48.570 4.280 ;
        RECT 49.410 0.835 49.950 4.280 ;
        RECT 50.790 0.835 51.790 4.280 ;
        RECT 52.630 0.835 53.170 4.280 ;
        RECT 54.010 0.835 55.010 4.280 ;
        RECT 55.850 0.835 56.390 4.280 ;
        RECT 57.230 0.835 58.230 4.280 ;
        RECT 59.070 0.835 59.610 4.280 ;
        RECT 60.450 0.835 61.450 4.280 ;
        RECT 62.290 0.835 62.830 4.280 ;
        RECT 63.670 0.835 64.670 4.280 ;
        RECT 65.510 0.835 66.050 4.280 ;
        RECT 66.890 0.835 67.890 4.280 ;
        RECT 68.730 0.835 69.270 4.280 ;
        RECT 70.110 0.835 71.110 4.280 ;
        RECT 71.950 0.835 72.490 4.280 ;
        RECT 73.330 0.835 74.330 4.280 ;
        RECT 75.170 0.835 75.710 4.280 ;
        RECT 76.550 0.835 77.550 4.280 ;
        RECT 78.390 0.835 78.930 4.280 ;
        RECT 79.770 0.835 80.770 4.280 ;
        RECT 81.610 0.835 82.150 4.280 ;
        RECT 82.990 0.835 83.990 4.280 ;
        RECT 84.830 0.835 85.370 4.280 ;
        RECT 86.210 0.835 87.210 4.280 ;
        RECT 88.050 0.835 88.590 4.280 ;
        RECT 89.430 0.835 90.430 4.280 ;
        RECT 91.270 0.835 91.810 4.280 ;
        RECT 92.650 0.835 93.650 4.280 ;
        RECT 94.490 0.835 95.030 4.280 ;
        RECT 95.870 0.835 96.870 4.280 ;
        RECT 97.710 0.835 98.250 4.280 ;
        RECT 99.090 0.835 100.090 4.280 ;
        RECT 100.930 0.835 101.930 4.280 ;
        RECT 102.770 0.835 103.310 4.280 ;
        RECT 104.150 0.835 105.150 4.280 ;
        RECT 105.990 0.835 106.530 4.280 ;
        RECT 107.370 0.835 108.370 4.280 ;
        RECT 109.210 0.835 109.750 4.280 ;
        RECT 110.590 0.835 111.590 4.280 ;
        RECT 112.430 0.835 112.970 4.280 ;
        RECT 113.810 0.835 114.810 4.280 ;
        RECT 115.650 0.835 116.190 4.280 ;
        RECT 117.030 0.835 118.030 4.280 ;
        RECT 118.870 0.835 119.410 4.280 ;
        RECT 120.250 0.835 121.250 4.280 ;
        RECT 122.090 0.835 122.630 4.280 ;
        RECT 123.470 0.835 124.470 4.280 ;
        RECT 125.310 0.835 125.850 4.280 ;
        RECT 126.690 0.835 127.690 4.280 ;
        RECT 128.530 0.835 129.070 4.280 ;
        RECT 129.910 0.835 130.910 4.280 ;
        RECT 131.750 0.835 132.290 4.280 ;
        RECT 133.130 0.835 134.130 4.280 ;
        RECT 134.970 0.835 135.510 4.280 ;
        RECT 136.350 0.835 137.350 4.280 ;
        RECT 138.190 0.835 138.730 4.280 ;
        RECT 139.570 0.835 140.570 4.280 ;
        RECT 141.410 0.835 141.950 4.280 ;
        RECT 142.790 0.835 143.790 4.280 ;
        RECT 144.630 0.835 145.170 4.280 ;
        RECT 146.010 0.835 147.010 4.280 ;
        RECT 147.850 0.835 148.390 4.280 ;
        RECT 149.230 0.835 150.230 4.280 ;
        RECT 151.070 0.835 151.610 4.280 ;
        RECT 152.450 0.835 153.450 4.280 ;
        RECT 154.290 0.835 154.830 4.280 ;
        RECT 155.670 0.835 156.670 4.280 ;
        RECT 157.510 0.835 158.050 4.280 ;
        RECT 158.890 0.835 159.890 4.280 ;
        RECT 160.730 0.835 161.270 4.280 ;
        RECT 162.110 0.835 163.110 4.280 ;
        RECT 163.950 0.835 164.490 4.280 ;
        RECT 165.330 0.835 166.330 4.280 ;
        RECT 167.170 0.835 167.710 4.280 ;
        RECT 168.550 0.835 169.550 4.280 ;
        RECT 170.390 0.835 170.930 4.280 ;
        RECT 171.770 0.835 172.770 4.280 ;
        RECT 173.610 0.835 174.150 4.280 ;
        RECT 174.990 0.835 175.990 4.280 ;
        RECT 176.830 0.835 177.370 4.280 ;
        RECT 178.210 0.835 179.210 4.280 ;
        RECT 180.050 0.835 180.590 4.280 ;
        RECT 181.430 0.835 182.430 4.280 ;
        RECT 183.270 0.835 183.810 4.280 ;
        RECT 184.650 0.835 185.650 4.280 ;
        RECT 186.490 0.835 187.030 4.280 ;
        RECT 187.870 0.835 188.870 4.280 ;
        RECT 189.710 0.835 190.250 4.280 ;
        RECT 191.090 0.835 192.090 4.280 ;
        RECT 192.930 0.835 193.470 4.280 ;
        RECT 194.310 0.835 195.310 4.280 ;
        RECT 196.150 0.835 196.690 4.280 ;
        RECT 197.530 0.835 198.530 4.280 ;
        RECT 199.370 0.835 200.370 4.280 ;
        RECT 201.210 0.835 201.750 4.280 ;
        RECT 202.590 0.835 203.590 4.280 ;
        RECT 204.430 0.835 204.970 4.280 ;
        RECT 205.810 0.835 206.810 4.280 ;
        RECT 207.650 0.835 208.190 4.280 ;
        RECT 209.030 0.835 210.030 4.280 ;
        RECT 210.870 0.835 211.410 4.280 ;
        RECT 212.250 0.835 213.250 4.280 ;
        RECT 214.090 0.835 214.630 4.280 ;
        RECT 215.470 0.835 216.470 4.280 ;
        RECT 217.310 0.835 217.850 4.280 ;
        RECT 218.690 0.835 219.690 4.280 ;
        RECT 220.530 0.835 221.070 4.280 ;
        RECT 221.910 0.835 222.910 4.280 ;
        RECT 223.750 0.835 224.290 4.280 ;
        RECT 225.130 0.835 226.130 4.280 ;
        RECT 226.970 0.835 227.510 4.280 ;
        RECT 228.350 0.835 229.350 4.280 ;
        RECT 230.190 0.835 230.730 4.280 ;
        RECT 231.570 0.835 232.570 4.280 ;
        RECT 233.410 0.835 233.950 4.280 ;
        RECT 234.790 0.835 235.790 4.280 ;
        RECT 236.630 0.835 237.170 4.280 ;
        RECT 238.010 0.835 239.010 4.280 ;
        RECT 239.850 0.835 240.390 4.280 ;
        RECT 241.230 0.835 242.230 4.280 ;
        RECT 243.070 0.835 243.610 4.280 ;
        RECT 244.450 0.835 245.450 4.280 ;
        RECT 246.290 0.835 246.830 4.280 ;
        RECT 247.670 0.835 248.670 4.280 ;
        RECT 249.510 0.835 250.050 4.280 ;
        RECT 250.890 0.835 251.890 4.280 ;
        RECT 252.730 0.835 253.270 4.280 ;
        RECT 254.110 0.835 255.110 4.280 ;
        RECT 255.950 0.835 256.490 4.280 ;
        RECT 257.330 0.835 258.330 4.280 ;
        RECT 259.170 0.835 259.710 4.280 ;
        RECT 260.550 0.835 261.550 4.280 ;
        RECT 262.390 0.835 262.930 4.280 ;
        RECT 263.770 0.835 264.770 4.280 ;
        RECT 265.610 0.835 266.150 4.280 ;
        RECT 266.990 0.835 267.990 4.280 ;
        RECT 268.830 0.835 269.370 4.280 ;
        RECT 270.210 0.835 271.210 4.280 ;
        RECT 272.050 0.835 272.590 4.280 ;
        RECT 273.430 0.835 274.430 4.280 ;
        RECT 275.270 0.835 275.810 4.280 ;
        RECT 276.650 0.835 277.650 4.280 ;
        RECT 278.490 0.835 279.030 4.280 ;
        RECT 279.870 0.835 280.870 4.280 ;
        RECT 281.710 0.835 282.250 4.280 ;
        RECT 283.090 0.835 284.090 4.280 ;
        RECT 284.930 0.835 285.470 4.280 ;
        RECT 286.310 0.835 287.310 4.280 ;
        RECT 288.150 0.835 288.690 4.280 ;
        RECT 289.530 0.835 290.530 4.280 ;
        RECT 291.370 0.835 291.910 4.280 ;
        RECT 292.750 0.835 293.750 4.280 ;
        RECT 294.590 0.835 295.130 4.280 ;
        RECT 295.970 0.835 296.970 4.280 ;
        RECT 297.810 0.835 298.350 4.280 ;
        RECT 299.190 0.835 300.190 4.280 ;
        RECT 301.030 0.835 302.030 4.280 ;
        RECT 302.870 0.835 303.410 4.280 ;
        RECT 304.250 0.835 305.250 4.280 ;
        RECT 306.090 0.835 306.630 4.280 ;
        RECT 307.470 0.835 308.470 4.280 ;
        RECT 309.310 0.835 309.850 4.280 ;
        RECT 310.690 0.835 311.690 4.280 ;
        RECT 312.530 0.835 313.070 4.280 ;
        RECT 313.910 0.835 314.910 4.280 ;
        RECT 315.750 0.835 316.290 4.280 ;
        RECT 317.130 0.835 318.130 4.280 ;
        RECT 318.970 0.835 319.510 4.280 ;
        RECT 320.350 0.835 321.350 4.280 ;
        RECT 322.190 0.835 322.730 4.280 ;
        RECT 323.570 0.835 324.570 4.280 ;
        RECT 325.410 0.835 325.950 4.280 ;
        RECT 326.790 0.835 327.790 4.280 ;
        RECT 328.630 0.835 329.170 4.280 ;
        RECT 330.010 0.835 331.010 4.280 ;
        RECT 331.850 0.835 332.390 4.280 ;
        RECT 333.230 0.835 334.230 4.280 ;
        RECT 335.070 0.835 335.610 4.280 ;
        RECT 336.450 0.835 337.450 4.280 ;
        RECT 338.290 0.835 338.830 4.280 ;
        RECT 339.670 0.835 340.670 4.280 ;
        RECT 341.510 0.835 342.050 4.280 ;
        RECT 342.890 0.835 343.890 4.280 ;
        RECT 344.730 0.835 345.270 4.280 ;
        RECT 346.110 0.835 347.110 4.280 ;
        RECT 347.950 0.835 348.490 4.280 ;
        RECT 349.330 0.835 350.330 4.280 ;
        RECT 351.170 0.835 351.710 4.280 ;
        RECT 352.550 0.835 353.550 4.280 ;
        RECT 354.390 0.835 354.930 4.280 ;
        RECT 355.770 0.835 356.770 4.280 ;
        RECT 357.610 0.835 358.150 4.280 ;
        RECT 358.990 0.835 359.990 4.280 ;
        RECT 360.830 0.835 361.370 4.280 ;
        RECT 362.210 0.835 363.210 4.280 ;
        RECT 364.050 0.835 364.590 4.280 ;
        RECT 365.430 0.835 366.430 4.280 ;
        RECT 367.270 0.835 367.810 4.280 ;
        RECT 368.650 0.835 369.650 4.280 ;
        RECT 370.490 0.835 371.030 4.280 ;
        RECT 371.870 0.835 372.870 4.280 ;
        RECT 373.710 0.835 374.250 4.280 ;
        RECT 375.090 0.835 376.090 4.280 ;
        RECT 376.930 0.835 377.470 4.280 ;
        RECT 378.310 0.835 379.310 4.280 ;
        RECT 380.150 0.835 380.690 4.280 ;
        RECT 381.530 0.835 382.530 4.280 ;
        RECT 383.370 0.835 383.910 4.280 ;
        RECT 384.750 0.835 385.750 4.280 ;
        RECT 386.590 0.835 387.130 4.280 ;
        RECT 387.970 0.835 388.970 4.280 ;
        RECT 389.810 0.835 390.350 4.280 ;
        RECT 391.190 0.835 392.190 4.280 ;
        RECT 393.030 0.835 393.570 4.280 ;
        RECT 394.410 0.835 395.410 4.280 ;
        RECT 396.250 0.835 396.790 4.280 ;
        RECT 397.630 0.835 398.630 4.280 ;
      LAYER met3 ;
        RECT 4.400 398.120 395.600 398.985 ;
        RECT 4.000 397.480 396.000 398.120 ;
        RECT 4.400 396.080 395.600 397.480 ;
        RECT 4.400 395.440 396.000 396.080 ;
        RECT 4.400 394.720 395.600 395.440 ;
        RECT 4.000 394.080 395.600 394.720 ;
        RECT 4.400 392.680 395.600 394.080 ;
        RECT 4.400 392.040 396.000 392.680 ;
        RECT 4.400 391.320 395.600 392.040 ;
        RECT 4.000 390.680 395.600 391.320 ;
        RECT 4.400 390.640 395.600 390.680 ;
        RECT 4.400 390.000 396.000 390.640 ;
        RECT 4.400 389.280 395.600 390.000 ;
        RECT 4.000 388.640 395.600 389.280 ;
        RECT 4.400 387.240 395.600 388.640 ;
        RECT 4.400 386.600 396.000 387.240 ;
        RECT 4.400 385.880 395.600 386.600 ;
        RECT 4.000 385.240 395.600 385.880 ;
        RECT 4.400 385.200 395.600 385.240 ;
        RECT 4.400 384.560 396.000 385.200 ;
        RECT 4.400 382.480 395.600 384.560 ;
        RECT 4.000 381.840 395.600 382.480 ;
        RECT 4.400 381.800 395.600 381.840 ;
        RECT 4.400 381.160 396.000 381.800 ;
        RECT 4.400 379.760 395.600 381.160 ;
        RECT 4.400 379.120 396.000 379.760 ;
        RECT 4.400 379.080 395.600 379.120 ;
        RECT 4.000 378.440 395.600 379.080 ;
        RECT 4.400 377.720 395.600 378.440 ;
        RECT 4.400 377.080 396.000 377.720 ;
        RECT 4.400 377.040 395.600 377.080 ;
        RECT 4.000 376.400 395.600 377.040 ;
        RECT 4.400 374.320 395.600 376.400 ;
        RECT 4.400 373.680 396.000 374.320 ;
        RECT 4.400 373.640 395.600 373.680 ;
        RECT 4.000 373.000 395.600 373.640 ;
        RECT 4.400 372.280 395.600 373.000 ;
        RECT 4.400 371.640 396.000 372.280 ;
        RECT 4.400 370.240 395.600 371.640 ;
        RECT 4.000 369.600 395.600 370.240 ;
        RECT 4.400 368.880 395.600 369.600 ;
        RECT 4.400 368.240 396.000 368.880 ;
        RECT 4.400 366.840 395.600 368.240 ;
        RECT 4.000 366.200 396.000 366.840 ;
        RECT 4.400 364.800 395.600 366.200 ;
        RECT 4.000 364.160 395.600 364.800 ;
        RECT 4.400 363.440 395.600 364.160 ;
        RECT 4.400 362.800 396.000 363.440 ;
        RECT 4.400 361.400 395.600 362.800 ;
        RECT 4.000 360.760 396.000 361.400 ;
        RECT 4.400 359.360 395.600 360.760 ;
        RECT 4.400 358.720 396.000 359.360 ;
        RECT 4.400 358.000 395.600 358.720 ;
        RECT 4.000 357.360 395.600 358.000 ;
        RECT 4.400 355.960 395.600 357.360 ;
        RECT 4.000 355.320 396.000 355.960 ;
        RECT 4.400 353.920 395.600 355.320 ;
        RECT 4.400 353.280 396.000 353.920 ;
        RECT 4.400 352.560 395.600 353.280 ;
        RECT 4.000 351.920 395.600 352.560 ;
        RECT 4.400 350.520 395.600 351.920 ;
        RECT 4.400 349.880 396.000 350.520 ;
        RECT 4.400 349.160 395.600 349.880 ;
        RECT 4.000 348.520 395.600 349.160 ;
        RECT 4.400 348.480 395.600 348.520 ;
        RECT 4.400 347.840 396.000 348.480 ;
        RECT 4.400 345.760 395.600 347.840 ;
        RECT 4.000 345.120 395.600 345.760 ;
        RECT 4.400 345.080 395.600 345.120 ;
        RECT 4.400 344.440 396.000 345.080 ;
        RECT 4.400 343.720 395.600 344.440 ;
        RECT 4.000 343.080 395.600 343.720 ;
        RECT 4.400 343.040 395.600 343.080 ;
        RECT 4.400 342.400 396.000 343.040 ;
        RECT 4.400 341.000 395.600 342.400 ;
        RECT 4.400 340.360 396.000 341.000 ;
        RECT 4.400 340.320 395.600 340.360 ;
        RECT 4.000 339.680 395.600 340.320 ;
        RECT 4.400 337.600 395.600 339.680 ;
        RECT 4.400 336.960 396.000 337.600 ;
        RECT 4.400 336.920 395.600 336.960 ;
        RECT 4.000 336.280 395.600 336.920 ;
        RECT 4.400 335.560 395.600 336.280 ;
        RECT 4.400 334.920 396.000 335.560 ;
        RECT 4.400 333.520 395.600 334.920 ;
        RECT 4.000 332.880 395.600 333.520 ;
        RECT 4.400 332.160 395.600 332.880 ;
        RECT 4.400 331.520 396.000 332.160 ;
        RECT 4.400 331.480 395.600 331.520 ;
        RECT 4.000 330.840 395.600 331.480 ;
        RECT 4.400 330.120 395.600 330.840 ;
        RECT 4.400 329.480 396.000 330.120 ;
        RECT 4.400 328.080 395.600 329.480 ;
        RECT 4.000 327.440 395.600 328.080 ;
        RECT 4.400 326.720 395.600 327.440 ;
        RECT 4.400 326.080 396.000 326.720 ;
        RECT 4.400 324.680 395.600 326.080 ;
        RECT 4.000 324.040 396.000 324.680 ;
        RECT 4.400 322.640 395.600 324.040 ;
        RECT 4.000 322.000 395.600 322.640 ;
        RECT 4.400 321.280 395.600 322.000 ;
        RECT 4.400 320.640 396.000 321.280 ;
        RECT 4.400 319.240 395.600 320.640 ;
        RECT 4.000 318.600 396.000 319.240 ;
        RECT 4.400 317.200 395.600 318.600 ;
        RECT 4.400 316.560 396.000 317.200 ;
        RECT 4.400 315.840 395.600 316.560 ;
        RECT 4.000 315.200 395.600 315.840 ;
        RECT 4.400 313.800 395.600 315.200 ;
        RECT 4.400 313.160 396.000 313.800 ;
        RECT 4.400 312.440 395.600 313.160 ;
        RECT 4.000 311.800 395.600 312.440 ;
        RECT 4.400 311.760 395.600 311.800 ;
        RECT 4.400 311.120 396.000 311.760 ;
        RECT 4.400 310.400 395.600 311.120 ;
        RECT 4.000 309.760 395.600 310.400 ;
        RECT 4.400 308.360 395.600 309.760 ;
        RECT 4.400 307.720 396.000 308.360 ;
        RECT 4.400 307.000 395.600 307.720 ;
        RECT 4.000 306.360 395.600 307.000 ;
        RECT 4.400 306.320 395.600 306.360 ;
        RECT 4.400 305.680 396.000 306.320 ;
        RECT 4.400 303.600 395.600 305.680 ;
        RECT 4.000 302.960 395.600 303.600 ;
        RECT 4.400 302.920 395.600 302.960 ;
        RECT 4.400 302.280 396.000 302.920 ;
        RECT 4.400 300.880 395.600 302.280 ;
        RECT 4.400 300.240 396.000 300.880 ;
        RECT 4.400 300.200 395.600 300.240 ;
        RECT 4.000 299.560 395.600 300.200 ;
        RECT 4.400 298.840 395.600 299.560 ;
        RECT 4.400 298.200 396.000 298.840 ;
        RECT 4.400 298.160 395.600 298.200 ;
        RECT 4.000 297.520 395.600 298.160 ;
        RECT 4.400 295.440 395.600 297.520 ;
        RECT 4.400 294.800 396.000 295.440 ;
        RECT 4.400 294.760 395.600 294.800 ;
        RECT 4.000 294.120 395.600 294.760 ;
        RECT 4.400 293.400 395.600 294.120 ;
        RECT 4.400 292.760 396.000 293.400 ;
        RECT 4.400 291.360 395.600 292.760 ;
        RECT 4.000 290.720 395.600 291.360 ;
        RECT 4.400 290.000 395.600 290.720 ;
        RECT 4.400 289.360 396.000 290.000 ;
        RECT 4.400 289.320 395.600 289.360 ;
        RECT 4.000 288.680 395.600 289.320 ;
        RECT 4.400 287.960 395.600 288.680 ;
        RECT 4.400 287.320 396.000 287.960 ;
        RECT 4.400 285.920 395.600 287.320 ;
        RECT 4.000 285.280 395.600 285.920 ;
        RECT 4.400 284.560 395.600 285.280 ;
        RECT 4.400 283.920 396.000 284.560 ;
        RECT 4.400 282.520 395.600 283.920 ;
        RECT 4.000 281.880 396.000 282.520 ;
        RECT 4.400 280.480 395.600 281.880 ;
        RECT 4.400 279.840 396.000 280.480 ;
        RECT 4.400 279.120 395.600 279.840 ;
        RECT 4.000 278.480 395.600 279.120 ;
        RECT 4.400 277.080 395.600 278.480 ;
        RECT 4.000 276.440 396.000 277.080 ;
        RECT 4.400 275.040 395.600 276.440 ;
        RECT 4.400 274.400 396.000 275.040 ;
        RECT 4.400 273.680 395.600 274.400 ;
        RECT 4.000 273.040 395.600 273.680 ;
        RECT 4.400 271.640 395.600 273.040 ;
        RECT 4.400 271.000 396.000 271.640 ;
        RECT 4.400 270.280 395.600 271.000 ;
        RECT 4.000 269.640 395.600 270.280 ;
        RECT 4.400 269.600 395.600 269.640 ;
        RECT 4.400 268.960 396.000 269.600 ;
        RECT 4.400 266.880 395.600 268.960 ;
        RECT 4.000 266.240 395.600 266.880 ;
        RECT 4.400 266.200 395.600 266.240 ;
        RECT 4.400 265.560 396.000 266.200 ;
        RECT 4.400 264.840 395.600 265.560 ;
        RECT 4.000 264.200 395.600 264.840 ;
        RECT 4.400 264.160 395.600 264.200 ;
        RECT 4.400 263.520 396.000 264.160 ;
        RECT 4.400 261.440 395.600 263.520 ;
        RECT 4.000 260.800 395.600 261.440 ;
        RECT 4.400 260.760 395.600 260.800 ;
        RECT 4.400 260.120 396.000 260.760 ;
        RECT 4.400 258.720 395.600 260.120 ;
        RECT 4.400 258.080 396.000 258.720 ;
        RECT 4.400 258.040 395.600 258.080 ;
        RECT 4.000 257.400 395.600 258.040 ;
        RECT 4.400 256.680 395.600 257.400 ;
        RECT 4.400 256.040 396.000 256.680 ;
        RECT 4.400 256.000 395.600 256.040 ;
        RECT 4.000 255.360 395.600 256.000 ;
        RECT 4.400 253.280 395.600 255.360 ;
        RECT 4.400 252.640 396.000 253.280 ;
        RECT 4.400 252.600 395.600 252.640 ;
        RECT 4.000 251.960 395.600 252.600 ;
        RECT 4.400 251.240 395.600 251.960 ;
        RECT 4.400 250.600 396.000 251.240 ;
        RECT 4.400 249.200 395.600 250.600 ;
        RECT 4.000 248.560 395.600 249.200 ;
        RECT 4.400 247.840 395.600 248.560 ;
        RECT 4.400 247.200 396.000 247.840 ;
        RECT 4.400 245.800 395.600 247.200 ;
        RECT 4.000 245.160 396.000 245.800 ;
        RECT 4.400 243.760 395.600 245.160 ;
        RECT 4.000 243.120 395.600 243.760 ;
        RECT 4.400 242.400 395.600 243.120 ;
        RECT 4.400 241.760 396.000 242.400 ;
        RECT 4.400 240.360 395.600 241.760 ;
        RECT 4.000 239.720 396.000 240.360 ;
        RECT 4.400 238.320 395.600 239.720 ;
        RECT 4.400 237.680 396.000 238.320 ;
        RECT 4.400 236.960 395.600 237.680 ;
        RECT 4.000 236.320 395.600 236.960 ;
        RECT 4.400 234.920 395.600 236.320 ;
        RECT 4.400 234.280 396.000 234.920 ;
        RECT 4.400 233.560 395.600 234.280 ;
        RECT 4.000 232.920 395.600 233.560 ;
        RECT 4.400 232.880 395.600 232.920 ;
        RECT 4.400 232.240 396.000 232.880 ;
        RECT 4.400 231.520 395.600 232.240 ;
        RECT 4.000 230.880 395.600 231.520 ;
        RECT 4.400 229.480 395.600 230.880 ;
        RECT 4.400 228.840 396.000 229.480 ;
        RECT 4.400 228.120 395.600 228.840 ;
        RECT 4.000 227.480 395.600 228.120 ;
        RECT 4.400 227.440 395.600 227.480 ;
        RECT 4.400 226.800 396.000 227.440 ;
        RECT 4.400 224.720 395.600 226.800 ;
        RECT 4.000 224.080 395.600 224.720 ;
        RECT 4.400 224.040 395.600 224.080 ;
        RECT 4.400 223.400 396.000 224.040 ;
        RECT 4.400 222.680 395.600 223.400 ;
        RECT 4.000 222.040 395.600 222.680 ;
        RECT 4.400 222.000 395.600 222.040 ;
        RECT 4.400 221.360 396.000 222.000 ;
        RECT 4.400 219.960 395.600 221.360 ;
        RECT 4.400 219.320 396.000 219.960 ;
        RECT 4.400 219.280 395.600 219.320 ;
        RECT 4.000 218.640 395.600 219.280 ;
        RECT 4.400 216.560 395.600 218.640 ;
        RECT 4.400 215.920 396.000 216.560 ;
        RECT 4.400 215.880 395.600 215.920 ;
        RECT 4.000 215.240 395.600 215.880 ;
        RECT 4.400 214.520 395.600 215.240 ;
        RECT 4.400 213.880 396.000 214.520 ;
        RECT 4.400 212.480 395.600 213.880 ;
        RECT 4.000 211.840 395.600 212.480 ;
        RECT 4.400 211.120 395.600 211.840 ;
        RECT 4.400 210.480 396.000 211.120 ;
        RECT 4.400 210.440 395.600 210.480 ;
        RECT 4.000 209.800 395.600 210.440 ;
        RECT 4.400 209.080 395.600 209.800 ;
        RECT 4.400 208.440 396.000 209.080 ;
        RECT 4.400 207.040 395.600 208.440 ;
        RECT 4.000 206.400 395.600 207.040 ;
        RECT 4.400 205.680 395.600 206.400 ;
        RECT 4.400 205.040 396.000 205.680 ;
        RECT 4.400 203.640 395.600 205.040 ;
        RECT 4.000 203.000 396.000 203.640 ;
        RECT 4.400 200.240 395.600 203.000 ;
        RECT 4.000 199.600 396.000 200.240 ;
        RECT 4.400 198.200 395.600 199.600 ;
        RECT 4.000 197.560 396.000 198.200 ;
        RECT 4.400 196.160 395.600 197.560 ;
        RECT 4.400 195.520 396.000 196.160 ;
        RECT 4.400 194.800 395.600 195.520 ;
        RECT 4.000 194.160 395.600 194.800 ;
        RECT 4.400 192.760 395.600 194.160 ;
        RECT 4.400 192.120 396.000 192.760 ;
        RECT 4.400 191.400 395.600 192.120 ;
        RECT 4.000 190.760 395.600 191.400 ;
        RECT 4.400 190.720 395.600 190.760 ;
        RECT 4.400 190.080 396.000 190.720 ;
        RECT 4.400 189.360 395.600 190.080 ;
        RECT 4.000 188.720 395.600 189.360 ;
        RECT 4.400 187.320 395.600 188.720 ;
        RECT 4.400 186.680 396.000 187.320 ;
        RECT 4.400 185.960 395.600 186.680 ;
        RECT 4.000 185.320 395.600 185.960 ;
        RECT 4.400 185.280 395.600 185.320 ;
        RECT 4.400 184.640 396.000 185.280 ;
        RECT 4.400 182.560 395.600 184.640 ;
        RECT 4.000 181.920 395.600 182.560 ;
        RECT 4.400 181.880 395.600 181.920 ;
        RECT 4.400 181.240 396.000 181.880 ;
        RECT 4.400 179.840 395.600 181.240 ;
        RECT 4.400 179.200 396.000 179.840 ;
        RECT 4.400 179.160 395.600 179.200 ;
        RECT 4.000 178.520 395.600 179.160 ;
        RECT 4.400 177.800 395.600 178.520 ;
        RECT 4.400 177.160 396.000 177.800 ;
        RECT 4.400 177.120 395.600 177.160 ;
        RECT 4.000 176.480 395.600 177.120 ;
        RECT 4.400 174.400 395.600 176.480 ;
        RECT 4.400 173.760 396.000 174.400 ;
        RECT 4.400 173.720 395.600 173.760 ;
        RECT 4.000 173.080 395.600 173.720 ;
        RECT 4.400 172.360 395.600 173.080 ;
        RECT 4.400 171.720 396.000 172.360 ;
        RECT 4.400 170.320 395.600 171.720 ;
        RECT 4.000 169.680 395.600 170.320 ;
        RECT 4.400 168.960 395.600 169.680 ;
        RECT 4.400 168.320 396.000 168.960 ;
        RECT 4.400 166.920 395.600 168.320 ;
        RECT 4.000 166.280 396.000 166.920 ;
        RECT 4.400 164.880 395.600 166.280 ;
        RECT 4.000 164.240 395.600 164.880 ;
        RECT 4.400 163.520 395.600 164.240 ;
        RECT 4.400 162.880 396.000 163.520 ;
        RECT 4.400 161.480 395.600 162.880 ;
        RECT 4.000 160.840 396.000 161.480 ;
        RECT 4.400 159.440 395.600 160.840 ;
        RECT 4.400 158.800 396.000 159.440 ;
        RECT 4.400 158.080 395.600 158.800 ;
        RECT 4.000 157.440 395.600 158.080 ;
        RECT 4.400 156.040 395.600 157.440 ;
        RECT 4.000 155.400 396.000 156.040 ;
        RECT 4.400 154.000 395.600 155.400 ;
        RECT 4.400 153.360 396.000 154.000 ;
        RECT 4.400 152.640 395.600 153.360 ;
        RECT 4.000 152.000 395.600 152.640 ;
        RECT 4.400 150.600 395.600 152.000 ;
        RECT 4.400 149.960 396.000 150.600 ;
        RECT 4.400 149.240 395.600 149.960 ;
        RECT 4.000 148.600 395.600 149.240 ;
        RECT 4.400 148.560 395.600 148.600 ;
        RECT 4.400 147.920 396.000 148.560 ;
        RECT 4.400 145.840 395.600 147.920 ;
        RECT 4.000 145.200 395.600 145.840 ;
        RECT 4.400 145.160 395.600 145.200 ;
        RECT 4.400 144.520 396.000 145.160 ;
        RECT 4.400 143.800 395.600 144.520 ;
        RECT 4.000 143.160 395.600 143.800 ;
        RECT 4.400 143.120 395.600 143.160 ;
        RECT 4.400 142.480 396.000 143.120 ;
        RECT 4.400 141.080 395.600 142.480 ;
        RECT 4.400 140.440 396.000 141.080 ;
        RECT 4.400 140.400 395.600 140.440 ;
        RECT 4.000 139.760 395.600 140.400 ;
        RECT 4.400 137.680 395.600 139.760 ;
        RECT 4.400 137.040 396.000 137.680 ;
        RECT 4.400 137.000 395.600 137.040 ;
        RECT 4.000 136.360 395.600 137.000 ;
        RECT 4.400 135.640 395.600 136.360 ;
        RECT 4.400 135.000 396.000 135.640 ;
        RECT 4.400 133.600 395.600 135.000 ;
        RECT 4.000 132.960 395.600 133.600 ;
        RECT 4.400 132.240 395.600 132.960 ;
        RECT 4.400 131.600 396.000 132.240 ;
        RECT 4.400 131.560 395.600 131.600 ;
        RECT 4.000 130.920 395.600 131.560 ;
        RECT 4.400 130.200 395.600 130.920 ;
        RECT 4.400 129.560 396.000 130.200 ;
        RECT 4.400 128.160 395.600 129.560 ;
        RECT 4.000 127.520 395.600 128.160 ;
        RECT 4.400 126.800 395.600 127.520 ;
        RECT 4.400 126.160 396.000 126.800 ;
        RECT 4.400 124.760 395.600 126.160 ;
        RECT 4.000 124.120 396.000 124.760 ;
        RECT 4.400 122.720 395.600 124.120 ;
        RECT 4.000 122.080 395.600 122.720 ;
        RECT 4.400 121.360 395.600 122.080 ;
        RECT 4.400 120.720 396.000 121.360 ;
        RECT 4.400 119.320 395.600 120.720 ;
        RECT 4.000 118.680 396.000 119.320 ;
        RECT 4.400 117.280 395.600 118.680 ;
        RECT 4.400 116.640 396.000 117.280 ;
        RECT 4.400 115.920 395.600 116.640 ;
        RECT 4.000 115.280 395.600 115.920 ;
        RECT 4.400 113.880 395.600 115.280 ;
        RECT 4.400 113.240 396.000 113.880 ;
        RECT 4.400 112.520 395.600 113.240 ;
        RECT 4.000 111.880 395.600 112.520 ;
        RECT 4.400 111.840 395.600 111.880 ;
        RECT 4.400 111.200 396.000 111.840 ;
        RECT 4.400 110.480 395.600 111.200 ;
        RECT 4.000 109.840 395.600 110.480 ;
        RECT 4.400 108.440 395.600 109.840 ;
        RECT 4.400 107.800 396.000 108.440 ;
        RECT 4.400 107.080 395.600 107.800 ;
        RECT 4.000 106.440 395.600 107.080 ;
        RECT 4.400 106.400 395.600 106.440 ;
        RECT 4.400 105.760 396.000 106.400 ;
        RECT 4.400 103.680 395.600 105.760 ;
        RECT 4.000 103.040 395.600 103.680 ;
        RECT 4.400 103.000 395.600 103.040 ;
        RECT 4.400 102.360 396.000 103.000 ;
        RECT 4.400 100.960 395.600 102.360 ;
        RECT 4.400 100.320 396.000 100.960 ;
        RECT 4.400 100.280 395.600 100.320 ;
        RECT 4.000 99.640 395.600 100.280 ;
        RECT 4.400 98.920 395.600 99.640 ;
        RECT 4.400 98.280 396.000 98.920 ;
        RECT 4.400 98.240 395.600 98.280 ;
        RECT 4.000 97.600 395.600 98.240 ;
        RECT 4.400 95.520 395.600 97.600 ;
        RECT 4.400 94.880 396.000 95.520 ;
        RECT 4.400 94.840 395.600 94.880 ;
        RECT 4.000 94.200 395.600 94.840 ;
        RECT 4.400 93.480 395.600 94.200 ;
        RECT 4.400 92.840 396.000 93.480 ;
        RECT 4.400 91.440 395.600 92.840 ;
        RECT 4.000 90.800 395.600 91.440 ;
        RECT 4.400 90.080 395.600 90.800 ;
        RECT 4.400 89.440 396.000 90.080 ;
        RECT 4.400 89.400 395.600 89.440 ;
        RECT 4.000 88.760 395.600 89.400 ;
        RECT 4.400 88.040 395.600 88.760 ;
        RECT 4.400 87.400 396.000 88.040 ;
        RECT 4.400 86.000 395.600 87.400 ;
        RECT 4.000 85.360 395.600 86.000 ;
        RECT 4.400 84.640 395.600 85.360 ;
        RECT 4.400 84.000 396.000 84.640 ;
        RECT 4.400 82.600 395.600 84.000 ;
        RECT 4.000 81.960 396.000 82.600 ;
        RECT 4.400 80.560 395.600 81.960 ;
        RECT 4.400 79.920 396.000 80.560 ;
        RECT 4.400 79.200 395.600 79.920 ;
        RECT 4.000 78.560 395.600 79.200 ;
        RECT 4.400 77.160 395.600 78.560 ;
        RECT 4.000 76.520 396.000 77.160 ;
        RECT 4.400 75.120 395.600 76.520 ;
        RECT 4.400 74.480 396.000 75.120 ;
        RECT 4.400 73.760 395.600 74.480 ;
        RECT 4.000 73.120 395.600 73.760 ;
        RECT 4.400 71.720 395.600 73.120 ;
        RECT 4.400 71.080 396.000 71.720 ;
        RECT 4.400 70.360 395.600 71.080 ;
        RECT 4.000 69.720 395.600 70.360 ;
        RECT 4.400 69.680 395.600 69.720 ;
        RECT 4.400 69.040 396.000 69.680 ;
        RECT 4.400 66.960 395.600 69.040 ;
        RECT 4.000 66.320 395.600 66.960 ;
        RECT 4.400 66.280 395.600 66.320 ;
        RECT 4.400 65.640 396.000 66.280 ;
        RECT 4.400 64.920 395.600 65.640 ;
        RECT 4.000 64.280 395.600 64.920 ;
        RECT 4.400 64.240 395.600 64.280 ;
        RECT 4.400 63.600 396.000 64.240 ;
        RECT 4.400 61.520 395.600 63.600 ;
        RECT 4.000 60.880 395.600 61.520 ;
        RECT 4.400 60.840 395.600 60.880 ;
        RECT 4.400 60.200 396.000 60.840 ;
        RECT 4.400 58.800 395.600 60.200 ;
        RECT 4.400 58.160 396.000 58.800 ;
        RECT 4.400 58.120 395.600 58.160 ;
        RECT 4.000 57.480 395.600 58.120 ;
        RECT 4.400 56.760 395.600 57.480 ;
        RECT 4.400 56.120 396.000 56.760 ;
        RECT 4.400 56.080 395.600 56.120 ;
        RECT 4.000 55.440 395.600 56.080 ;
        RECT 4.400 53.360 395.600 55.440 ;
        RECT 4.400 52.720 396.000 53.360 ;
        RECT 4.400 52.680 395.600 52.720 ;
        RECT 4.000 52.040 395.600 52.680 ;
        RECT 4.400 51.320 395.600 52.040 ;
        RECT 4.400 50.680 396.000 51.320 ;
        RECT 4.400 49.280 395.600 50.680 ;
        RECT 4.000 48.640 395.600 49.280 ;
        RECT 4.400 47.920 395.600 48.640 ;
        RECT 4.400 47.280 396.000 47.920 ;
        RECT 4.400 45.880 395.600 47.280 ;
        RECT 4.000 45.240 396.000 45.880 ;
        RECT 4.400 43.840 395.600 45.240 ;
        RECT 4.000 43.200 395.600 43.840 ;
        RECT 4.400 42.480 395.600 43.200 ;
        RECT 4.400 41.840 396.000 42.480 ;
        RECT 4.400 40.440 395.600 41.840 ;
        RECT 4.000 39.800 396.000 40.440 ;
        RECT 4.400 38.400 395.600 39.800 ;
        RECT 4.400 37.760 396.000 38.400 ;
        RECT 4.400 37.040 395.600 37.760 ;
        RECT 4.000 36.400 395.600 37.040 ;
        RECT 4.400 35.000 395.600 36.400 ;
        RECT 4.400 34.360 396.000 35.000 ;
        RECT 4.400 33.640 395.600 34.360 ;
        RECT 4.000 33.000 395.600 33.640 ;
        RECT 4.400 32.960 395.600 33.000 ;
        RECT 4.400 32.320 396.000 32.960 ;
        RECT 4.400 31.600 395.600 32.320 ;
        RECT 4.000 30.960 395.600 31.600 ;
        RECT 4.400 29.560 395.600 30.960 ;
        RECT 4.400 28.920 396.000 29.560 ;
        RECT 4.400 28.200 395.600 28.920 ;
        RECT 4.000 27.560 395.600 28.200 ;
        RECT 4.400 27.520 395.600 27.560 ;
        RECT 4.400 26.880 396.000 27.520 ;
        RECT 4.400 24.800 395.600 26.880 ;
        RECT 4.000 24.160 395.600 24.800 ;
        RECT 4.400 24.120 395.600 24.160 ;
        RECT 4.400 23.480 396.000 24.120 ;
        RECT 4.400 22.760 395.600 23.480 ;
        RECT 4.000 22.120 395.600 22.760 ;
        RECT 4.400 22.080 395.600 22.120 ;
        RECT 4.400 21.440 396.000 22.080 ;
        RECT 4.400 20.040 395.600 21.440 ;
        RECT 4.400 19.400 396.000 20.040 ;
        RECT 4.400 19.360 395.600 19.400 ;
        RECT 4.000 18.720 395.600 19.360 ;
        RECT 4.400 16.640 395.600 18.720 ;
        RECT 4.400 16.000 396.000 16.640 ;
        RECT 4.400 15.960 395.600 16.000 ;
        RECT 4.000 15.320 395.600 15.960 ;
        RECT 4.400 14.600 395.600 15.320 ;
        RECT 4.400 13.960 396.000 14.600 ;
        RECT 4.400 12.560 395.600 13.960 ;
        RECT 4.000 11.920 395.600 12.560 ;
        RECT 4.400 11.200 395.600 11.920 ;
        RECT 4.400 10.560 396.000 11.200 ;
        RECT 4.400 10.520 395.600 10.560 ;
        RECT 4.000 9.880 395.600 10.520 ;
        RECT 4.400 9.160 395.600 9.880 ;
        RECT 4.400 8.520 396.000 9.160 ;
        RECT 4.400 7.120 395.600 8.520 ;
        RECT 4.000 6.480 395.600 7.120 ;
        RECT 4.400 5.760 395.600 6.480 ;
        RECT 4.400 5.120 396.000 5.760 ;
        RECT 4.400 3.720 395.600 5.120 ;
        RECT 4.000 3.080 396.000 3.720 ;
        RECT 4.400 0.855 395.600 3.080 ;
      LAYER met4 ;
        RECT 8.575 11.735 20.640 364.985 ;
        RECT 23.040 11.735 97.440 364.985 ;
        RECT 99.840 11.735 174.240 364.985 ;
        RECT 176.640 11.735 251.040 364.985 ;
        RECT 253.440 11.735 323.545 364.985 ;
  END
END chip_controller
END LIBRARY

