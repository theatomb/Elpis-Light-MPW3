VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO custom_sram
  CLASS BLOCK ;
  FOREIGN custom_sram ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1500.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1263.480 4.000 1264.080 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 1496.000 595.610 1500.000 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 1496.000 243.250 1500.000 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 160.520 1200.000 161.120 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1202.280 1200.000 1202.880 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 235.320 1200.000 235.920 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1350.520 1200.000 1351.120 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1487.880 4.000 1488.480 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1052.680 1200.000 1053.280 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 904.440 1200.000 905.040 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.170 1496.000 1149.450 1500.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 458.360 1200.000 458.960 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 1496.000 545.010 1500.000 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END a[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.970 0.000 956.250 4.000 ;
    END
  END clk
  PIN csb0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.570 0.000 1006.850 4.000 ;
    END
  END csb0_to_sram
  PIN d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 1496.000 797.090 1500.000 ;
    END
  END d[0]
  PIN d[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 979.240 1200.000 979.840 ;
    END
  END d[10]
  PIN d[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END d[11]
  PIN d[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 967.000 4.000 967.600 ;
    END
  END d[12]
  PIN d[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 531.800 1200.000 532.400 ;
    END
  END d[13]
  PIN d[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 1496.000 695.890 1500.000 ;
    END
  END d[14]
  PIN d[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END d[15]
  PIN d[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 1496.000 897.370 1500.000 ;
    END
  END d[16]
  PIN d[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END d[17]
  PIN d[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1127.480 1200.000 1128.080 ;
    END
  END d[18]
  PIN d[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END d[19]
  PIN d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 1496.000 646.210 1500.000 ;
    END
  END d[1]
  PIN d[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END d[20]
  PIN d[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END d[21]
  PIN d[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 1496.000 847.690 1500.000 ;
    END
  END d[22]
  PIN d[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 1496.000 1048.250 1500.000 ;
    END
  END d[23]
  PIN d[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 1496.000 92.370 1500.000 ;
    END
  END d[24]
  PIN d[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 1496.000 142.970 1500.000 ;
    END
  END d[25]
  PIN d[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END d[26]
  PIN d[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END d[27]
  PIN d[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1275.720 1200.000 1276.320 ;
    END
  END d[28]
  PIN d[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END d[29]
  PIN d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END d[2]
  PIN d[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END d[30]
  PIN d[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 0.000 905.650 4.000 ;
    END
  END d[31]
  PIN d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 383.560 1200.000 384.160 ;
    END
  END d[3]
  PIN d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 85.720 1200.000 86.320 ;
    END
  END d[4]
  PIN d[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END d[5]
  PIN d[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 1496.000 41.770 1500.000 ;
    END
  END d[6]
  PIN d[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 0.000 1107.130 4.000 ;
    END
  END d[7]
  PIN d[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 1496.000 394.130 1500.000 ;
    END
  END d[8]
  PIN d[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 308.760 1200.000 309.360 ;
    END
  END d[9]
  PIN q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 681.400 1200.000 682.000 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END q[11]
  PIN q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 1496.000 293.850 1500.000 ;
    END
  END q[12]
  PIN q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 1496.000 495.330 1500.000 ;
    END
  END q[13]
  PIN q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1338.280 4.000 1338.880 ;
    END
  END q[14]
  PIN q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END q[15]
  PIN q[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END q[16]
  PIN q[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 1496.000 444.730 1500.000 ;
    END
  END q[17]
  PIN q[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 1496.000 746.490 1500.000 ;
    END
  END q[18]
  PIN q[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 1496.000 1098.850 1500.000 ;
    END
  END q[19]
  PIN q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END q[1]
  PIN q[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END q[20]
  PIN q[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END q[21]
  PIN q[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.850 1496.000 1199.130 1500.000 ;
    END
  END q[22]
  PIN q[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END q[23]
  PIN q[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END q[24]
  PIN q[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1425.320 1200.000 1425.920 ;
    END
  END q[25]
  PIN q[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 10.920 1200.000 11.520 ;
    END
  END q[26]
  PIN q[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END q[27]
  PIN q[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 754.840 1200.000 755.440 ;
    END
  END q[28]
  PIN q[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END q[29]
  PIN q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END q[2]
  PIN q[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END q[30]
  PIN q[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 829.640 1200.000 830.240 ;
    END
  END q[31]
  PIN q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 1496.000 998.570 1500.000 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.690 1496.000 947.970 1500.000 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 1496.000 192.650 1500.000 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 1496.000 344.450 1500.000 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END q[9]
  PIN spare_wen0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1413.080 4.000 1413.680 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
  END vssd1
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 606.600 1200.000 607.200 ;
    END
  END we
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.935 1487.925 ;
      LAYER met1 ;
        RECT 0.070 10.640 1199.150 1488.480 ;
      LAYER met2 ;
        RECT 0.100 1495.720 41.210 1496.000 ;
        RECT 42.050 1495.720 91.810 1496.000 ;
        RECT 92.650 1495.720 142.410 1496.000 ;
        RECT 143.250 1495.720 192.090 1496.000 ;
        RECT 192.930 1495.720 242.690 1496.000 ;
        RECT 243.530 1495.720 293.290 1496.000 ;
        RECT 294.130 1495.720 343.890 1496.000 ;
        RECT 344.730 1495.720 393.570 1496.000 ;
        RECT 394.410 1495.720 444.170 1496.000 ;
        RECT 445.010 1495.720 494.770 1496.000 ;
        RECT 495.610 1495.720 544.450 1496.000 ;
        RECT 545.290 1495.720 595.050 1496.000 ;
        RECT 595.890 1495.720 645.650 1496.000 ;
        RECT 646.490 1495.720 695.330 1496.000 ;
        RECT 696.170 1495.720 745.930 1496.000 ;
        RECT 746.770 1495.720 796.530 1496.000 ;
        RECT 797.370 1495.720 847.130 1496.000 ;
        RECT 847.970 1495.720 896.810 1496.000 ;
        RECT 897.650 1495.720 947.410 1496.000 ;
        RECT 948.250 1495.720 998.010 1496.000 ;
        RECT 998.850 1495.720 1047.690 1496.000 ;
        RECT 1048.530 1495.720 1098.290 1496.000 ;
        RECT 1099.130 1495.720 1148.890 1496.000 ;
        RECT 1149.730 1495.720 1198.570 1496.000 ;
        RECT 0.100 4.280 1199.120 1495.720 ;
        RECT 0.650 3.670 49.490 4.280 ;
        RECT 50.330 3.670 100.090 4.280 ;
        RECT 100.930 3.670 150.690 4.280 ;
        RECT 151.530 3.670 200.370 4.280 ;
        RECT 201.210 3.670 250.970 4.280 ;
        RECT 251.810 3.670 301.570 4.280 ;
        RECT 302.410 3.670 351.250 4.280 ;
        RECT 352.090 3.670 401.850 4.280 ;
        RECT 402.690 3.670 452.450 4.280 ;
        RECT 453.290 3.670 503.050 4.280 ;
        RECT 503.890 3.670 552.730 4.280 ;
        RECT 553.570 3.670 603.330 4.280 ;
        RECT 604.170 3.670 653.930 4.280 ;
        RECT 654.770 3.670 703.610 4.280 ;
        RECT 704.450 3.670 754.210 4.280 ;
        RECT 755.050 3.670 804.810 4.280 ;
        RECT 805.650 3.670 854.490 4.280 ;
        RECT 855.330 3.670 905.090 4.280 ;
        RECT 905.930 3.670 955.690 4.280 ;
        RECT 956.530 3.670 1006.290 4.280 ;
        RECT 1007.130 3.670 1055.970 4.280 ;
        RECT 1056.810 3.670 1106.570 4.280 ;
        RECT 1107.410 3.670 1157.170 4.280 ;
        RECT 1158.010 3.670 1199.120 4.280 ;
      LAYER met3 ;
        RECT 4.400 1487.480 1196.000 1488.005 ;
        RECT 4.000 1426.320 1196.000 1487.480 ;
        RECT 4.000 1424.920 1195.600 1426.320 ;
        RECT 4.000 1414.080 1196.000 1424.920 ;
        RECT 4.400 1412.680 1196.000 1414.080 ;
        RECT 4.000 1351.520 1196.000 1412.680 ;
        RECT 4.000 1350.120 1195.600 1351.520 ;
        RECT 4.000 1339.280 1196.000 1350.120 ;
        RECT 4.400 1337.880 1196.000 1339.280 ;
        RECT 4.000 1276.720 1196.000 1337.880 ;
        RECT 4.000 1275.320 1195.600 1276.720 ;
        RECT 4.000 1264.480 1196.000 1275.320 ;
        RECT 4.400 1263.080 1196.000 1264.480 ;
        RECT 4.000 1203.280 1196.000 1263.080 ;
        RECT 4.000 1201.880 1195.600 1203.280 ;
        RECT 4.000 1191.040 1196.000 1201.880 ;
        RECT 4.400 1189.640 1196.000 1191.040 ;
        RECT 4.000 1128.480 1196.000 1189.640 ;
        RECT 4.000 1127.080 1195.600 1128.480 ;
        RECT 4.000 1116.240 1196.000 1127.080 ;
        RECT 4.400 1114.840 1196.000 1116.240 ;
        RECT 4.000 1053.680 1196.000 1114.840 ;
        RECT 4.000 1052.280 1195.600 1053.680 ;
        RECT 4.000 1041.440 1196.000 1052.280 ;
        RECT 4.400 1040.040 1196.000 1041.440 ;
        RECT 4.000 980.240 1196.000 1040.040 ;
        RECT 4.000 978.840 1195.600 980.240 ;
        RECT 4.000 968.000 1196.000 978.840 ;
        RECT 4.400 966.600 1196.000 968.000 ;
        RECT 4.000 905.440 1196.000 966.600 ;
        RECT 4.000 904.040 1195.600 905.440 ;
        RECT 4.000 893.200 1196.000 904.040 ;
        RECT 4.400 891.800 1196.000 893.200 ;
        RECT 4.000 830.640 1196.000 891.800 ;
        RECT 4.000 829.240 1195.600 830.640 ;
        RECT 4.000 818.400 1196.000 829.240 ;
        RECT 4.400 817.000 1196.000 818.400 ;
        RECT 4.000 755.840 1196.000 817.000 ;
        RECT 4.000 754.440 1195.600 755.840 ;
        RECT 4.000 744.960 1196.000 754.440 ;
        RECT 4.400 743.560 1196.000 744.960 ;
        RECT 4.000 682.400 1196.000 743.560 ;
        RECT 4.000 681.000 1195.600 682.400 ;
        RECT 4.000 670.160 1196.000 681.000 ;
        RECT 4.400 668.760 1196.000 670.160 ;
        RECT 4.000 607.600 1196.000 668.760 ;
        RECT 4.000 606.200 1195.600 607.600 ;
        RECT 4.000 595.360 1196.000 606.200 ;
        RECT 4.400 593.960 1196.000 595.360 ;
        RECT 4.000 532.800 1196.000 593.960 ;
        RECT 4.000 531.400 1195.600 532.800 ;
        RECT 4.000 520.560 1196.000 531.400 ;
        RECT 4.400 519.160 1196.000 520.560 ;
        RECT 4.000 459.360 1196.000 519.160 ;
        RECT 4.000 457.960 1195.600 459.360 ;
        RECT 4.000 447.120 1196.000 457.960 ;
        RECT 4.400 445.720 1196.000 447.120 ;
        RECT 4.000 384.560 1196.000 445.720 ;
        RECT 4.000 383.160 1195.600 384.560 ;
        RECT 4.000 372.320 1196.000 383.160 ;
        RECT 4.400 370.920 1196.000 372.320 ;
        RECT 4.000 309.760 1196.000 370.920 ;
        RECT 4.000 308.360 1195.600 309.760 ;
        RECT 4.000 297.520 1196.000 308.360 ;
        RECT 4.400 296.120 1196.000 297.520 ;
        RECT 4.000 236.320 1196.000 296.120 ;
        RECT 4.000 234.920 1195.600 236.320 ;
        RECT 4.000 224.080 1196.000 234.920 ;
        RECT 4.400 222.680 1196.000 224.080 ;
        RECT 4.000 161.520 1196.000 222.680 ;
        RECT 4.000 160.120 1195.600 161.520 ;
        RECT 4.000 149.280 1196.000 160.120 ;
        RECT 4.400 147.880 1196.000 149.280 ;
        RECT 4.000 86.720 1196.000 147.880 ;
        RECT 4.000 85.320 1195.600 86.720 ;
        RECT 4.000 74.480 1196.000 85.320 ;
        RECT 4.400 73.080 1196.000 74.480 ;
        RECT 4.000 11.920 1196.000 73.080 ;
        RECT 4.000 10.715 1195.600 11.920 ;
      LAYER met4 ;
        RECT 47.215 17.175 97.440 1480.865 ;
        RECT 99.840 17.175 174.240 1480.865 ;
        RECT 176.640 17.175 251.040 1480.865 ;
        RECT 253.440 17.175 327.840 1480.865 ;
        RECT 330.240 17.175 404.640 1480.865 ;
        RECT 407.040 17.175 481.440 1480.865 ;
        RECT 483.840 17.175 558.240 1480.865 ;
        RECT 560.640 17.175 635.040 1480.865 ;
        RECT 637.440 17.175 711.840 1480.865 ;
        RECT 714.240 17.175 788.640 1480.865 ;
        RECT 791.040 17.175 865.440 1480.865 ;
        RECT 867.840 17.175 942.240 1480.865 ;
        RECT 944.640 17.175 1019.040 1480.865 ;
        RECT 1021.440 17.175 1095.840 1480.865 ;
        RECT 1098.240 17.175 1113.825 1480.865 ;
  END
END custom_sram
END LIBRARY

