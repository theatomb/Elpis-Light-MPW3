VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO custom_sram
  CLASS BLOCK ;
  FOREIGN custom_sram ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1500.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 562.400 1200.000 563.000 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 862.280 1200.000 862.880 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 1496.000 599.750 1500.000 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 1496.000 670.590 1500.000 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1162.160 1200.000 1162.760 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 1496.000 811.810 1500.000 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 1496.000 176.090 1500.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 37.440 1200.000 38.040 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 187.040 1200.000 187.640 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END a[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END clk
  PIN csb0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END csb0_to_sram
  PIN d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END d[0]
  PIN d[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END d[10]
  PIN d[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 712.000 1200.000 712.600 ;
    END
  END d[11]
  PIN d[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 937.080 1200.000 937.680 ;
    END
  END d[12]
  PIN d[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END d[13]
  PIN d[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END d[14]
  PIN d[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END d[15]
  PIN d[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.760 4.000 904.360 ;
    END
  END d[16]
  PIN d[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1087.360 1200.000 1087.960 ;
    END
  END d[17]
  PIN d[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 1496.000 740.970 1500.000 ;
    END
  END d[18]
  PIN d[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END d[19]
  PIN d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 1496.000 105.710 1500.000 ;
    END
  END d[1]
  PIN d[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 0.000 882.190 4.000 ;
    END
  END d[20]
  PIN d[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1080.560 4.000 1081.160 ;
    END
  END d[21]
  PIN d[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.760 4.000 1125.360 ;
    END
  END d[22]
  PIN d[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 1496.000 953.030 1500.000 ;
    END
  END d[23]
  PIN d[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1212.480 4.000 1213.080 ;
    END
  END d[24]
  PIN d[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 1496.000 1023.410 1500.000 ;
    END
  END d[25]
  PIN d[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1345.080 4.000 1345.680 ;
    END
  END d[26]
  PIN d[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1389.280 4.000 1389.880 ;
    END
  END d[27]
  PIN d[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1433.480 4.000 1434.080 ;
    END
  END d[28]
  PIN d[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 1496.000 1094.250 1500.000 ;
    END
  END d[29]
  PIN d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END d[2]
  PIN d[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END d[30]
  PIN d[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1462.040 1200.000 1462.640 ;
    END
  END d[31]
  PIN d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END d[3]
  PIN d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END d[4]
  PIN d[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END d[5]
  PIN d[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 261.840 1200.000 262.440 ;
    END
  END d[6]
  PIN d[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 1496.000 317.310 1500.000 ;
    END
  END d[7]
  PIN d[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 412.120 1200.000 412.720 ;
    END
  END d[8]
  PIN d[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 1496.000 458.530 1500.000 ;
    END
  END d[9]
  PIN q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 1496.000 35.330 1500.000 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 637.200 1200.000 637.800 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 787.480 1200.000 788.080 ;
    END
  END q[11]
  PIN q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END q[12]
  PIN q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1011.880 1200.000 1012.480 ;
    END
  END q[13]
  PIN q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END q[14]
  PIN q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END q[15]
  PIN q[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END q[16]
  PIN q[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.160 4.000 992.760 ;
    END
  END q[17]
  PIN q[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END q[18]
  PIN q[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END q[19]
  PIN q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END q[1]
  PIN q[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 1496.000 882.190 1500.000 ;
    END
  END q[20]
  PIN q[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1236.960 1200.000 1237.560 ;
    END
  END q[21]
  PIN q[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1312.440 1200.000 1313.040 ;
    END
  END q[22]
  PIN q[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1168.280 4.000 1168.880 ;
    END
  END q[23]
  PIN q[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1256.680 4.000 1257.280 ;
    END
  END q[24]
  PIN q[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.880 4.000 1301.480 ;
    END
  END q[25]
  PIN q[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1387.240 1200.000 1387.840 ;
    END
  END q[26]
  PIN q[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.750 0.000 953.030 4.000 ;
    END
  END q[27]
  PIN q[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.130 0.000 1023.410 4.000 ;
    END
  END q[28]
  PIN q[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END q[29]
  PIN q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END q[2]
  PIN q[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 1496.000 1164.630 1500.000 ;
    END
  END q[30]
  PIN q[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1477.680 4.000 1478.280 ;
    END
  END q[31]
  PIN q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 1496.000 246.930 1500.000 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 112.240 1200.000 112.840 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 337.320 1200.000 337.920 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 1496.000 388.150 1500.000 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 486.920 1200.000 487.520 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 1496.000 529.370 1500.000 ;
    END
  END q[9]
  PIN spare_wen0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
  END vssd1
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END we
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1196.315 1487.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 1196.375 1488.080 ;
      LAYER met2 ;
        RECT 6.990 1495.720 34.770 1496.410 ;
        RECT 35.610 1495.720 105.150 1496.410 ;
        RECT 105.990 1495.720 175.530 1496.410 ;
        RECT 176.370 1495.720 246.370 1496.410 ;
        RECT 247.210 1495.720 316.750 1496.410 ;
        RECT 317.590 1495.720 387.590 1496.410 ;
        RECT 388.430 1495.720 457.970 1496.410 ;
        RECT 458.810 1495.720 528.810 1496.410 ;
        RECT 529.650 1495.720 599.190 1496.410 ;
        RECT 600.030 1495.720 670.030 1496.410 ;
        RECT 670.870 1495.720 740.410 1496.410 ;
        RECT 741.250 1495.720 811.250 1496.410 ;
        RECT 812.090 1495.720 881.630 1496.410 ;
        RECT 882.470 1495.720 952.470 1496.410 ;
        RECT 953.310 1495.720 1022.850 1496.410 ;
        RECT 1023.690 1495.720 1093.690 1496.410 ;
        RECT 1094.530 1495.720 1164.070 1496.410 ;
        RECT 1164.910 1495.720 1191.770 1496.410 ;
        RECT 6.990 4.280 1191.770 1495.720 ;
        RECT 6.990 4.000 34.770 4.280 ;
        RECT 35.610 4.000 105.150 4.280 ;
        RECT 105.990 4.000 175.530 4.280 ;
        RECT 176.370 4.000 246.370 4.280 ;
        RECT 247.210 4.000 316.750 4.280 ;
        RECT 317.590 4.000 387.590 4.280 ;
        RECT 388.430 4.000 457.970 4.280 ;
        RECT 458.810 4.000 528.810 4.280 ;
        RECT 529.650 4.000 599.190 4.280 ;
        RECT 600.030 4.000 670.030 4.280 ;
        RECT 670.870 4.000 740.410 4.280 ;
        RECT 741.250 4.000 811.250 4.280 ;
        RECT 812.090 4.000 881.630 4.280 ;
        RECT 882.470 4.000 952.470 4.280 ;
        RECT 953.310 4.000 1022.850 4.280 ;
        RECT 1023.690 4.000 1093.690 4.280 ;
        RECT 1094.530 4.000 1164.070 4.280 ;
        RECT 1164.910 4.000 1191.770 4.280 ;
      LAYER met3 ;
        RECT 4.000 1478.680 1196.000 1488.005 ;
        RECT 4.400 1477.280 1196.000 1478.680 ;
        RECT 4.000 1463.040 1196.000 1477.280 ;
        RECT 4.000 1461.640 1195.600 1463.040 ;
        RECT 4.000 1434.480 1196.000 1461.640 ;
        RECT 4.400 1433.080 1196.000 1434.480 ;
        RECT 4.000 1390.280 1196.000 1433.080 ;
        RECT 4.400 1388.880 1196.000 1390.280 ;
        RECT 4.000 1388.240 1196.000 1388.880 ;
        RECT 4.000 1386.840 1195.600 1388.240 ;
        RECT 4.000 1346.080 1196.000 1386.840 ;
        RECT 4.400 1344.680 1196.000 1346.080 ;
        RECT 4.000 1313.440 1196.000 1344.680 ;
        RECT 4.000 1312.040 1195.600 1313.440 ;
        RECT 4.000 1301.880 1196.000 1312.040 ;
        RECT 4.400 1300.480 1196.000 1301.880 ;
        RECT 4.000 1257.680 1196.000 1300.480 ;
        RECT 4.400 1256.280 1196.000 1257.680 ;
        RECT 4.000 1237.960 1196.000 1256.280 ;
        RECT 4.000 1236.560 1195.600 1237.960 ;
        RECT 4.000 1213.480 1196.000 1236.560 ;
        RECT 4.400 1212.080 1196.000 1213.480 ;
        RECT 4.000 1169.280 1196.000 1212.080 ;
        RECT 4.400 1167.880 1196.000 1169.280 ;
        RECT 4.000 1163.160 1196.000 1167.880 ;
        RECT 4.000 1161.760 1195.600 1163.160 ;
        RECT 4.000 1125.760 1196.000 1161.760 ;
        RECT 4.400 1124.360 1196.000 1125.760 ;
        RECT 4.000 1088.360 1196.000 1124.360 ;
        RECT 4.000 1086.960 1195.600 1088.360 ;
        RECT 4.000 1081.560 1196.000 1086.960 ;
        RECT 4.400 1080.160 1196.000 1081.560 ;
        RECT 4.000 1037.360 1196.000 1080.160 ;
        RECT 4.400 1035.960 1196.000 1037.360 ;
        RECT 4.000 1012.880 1196.000 1035.960 ;
        RECT 4.000 1011.480 1195.600 1012.880 ;
        RECT 4.000 993.160 1196.000 1011.480 ;
        RECT 4.400 991.760 1196.000 993.160 ;
        RECT 4.000 948.960 1196.000 991.760 ;
        RECT 4.400 947.560 1196.000 948.960 ;
        RECT 4.000 938.080 1196.000 947.560 ;
        RECT 4.000 936.680 1195.600 938.080 ;
        RECT 4.000 904.760 1196.000 936.680 ;
        RECT 4.400 903.360 1196.000 904.760 ;
        RECT 4.000 863.280 1196.000 903.360 ;
        RECT 4.000 861.880 1195.600 863.280 ;
        RECT 4.000 860.560 1196.000 861.880 ;
        RECT 4.400 859.160 1196.000 860.560 ;
        RECT 4.000 816.360 1196.000 859.160 ;
        RECT 4.400 814.960 1196.000 816.360 ;
        RECT 4.000 788.480 1196.000 814.960 ;
        RECT 4.000 787.080 1195.600 788.480 ;
        RECT 4.000 772.840 1196.000 787.080 ;
        RECT 4.400 771.440 1196.000 772.840 ;
        RECT 4.000 728.640 1196.000 771.440 ;
        RECT 4.400 727.240 1196.000 728.640 ;
        RECT 4.000 713.000 1196.000 727.240 ;
        RECT 4.000 711.600 1195.600 713.000 ;
        RECT 4.000 684.440 1196.000 711.600 ;
        RECT 4.400 683.040 1196.000 684.440 ;
        RECT 4.000 640.240 1196.000 683.040 ;
        RECT 4.400 638.840 1196.000 640.240 ;
        RECT 4.000 638.200 1196.000 638.840 ;
        RECT 4.000 636.800 1195.600 638.200 ;
        RECT 4.000 596.040 1196.000 636.800 ;
        RECT 4.400 594.640 1196.000 596.040 ;
        RECT 4.000 563.400 1196.000 594.640 ;
        RECT 4.000 562.000 1195.600 563.400 ;
        RECT 4.000 551.840 1196.000 562.000 ;
        RECT 4.400 550.440 1196.000 551.840 ;
        RECT 4.000 507.640 1196.000 550.440 ;
        RECT 4.400 506.240 1196.000 507.640 ;
        RECT 4.000 487.920 1196.000 506.240 ;
        RECT 4.000 486.520 1195.600 487.920 ;
        RECT 4.000 463.440 1196.000 486.520 ;
        RECT 4.400 462.040 1196.000 463.440 ;
        RECT 4.000 419.240 1196.000 462.040 ;
        RECT 4.400 417.840 1196.000 419.240 ;
        RECT 4.000 413.120 1196.000 417.840 ;
        RECT 4.000 411.720 1195.600 413.120 ;
        RECT 4.000 375.720 1196.000 411.720 ;
        RECT 4.400 374.320 1196.000 375.720 ;
        RECT 4.000 338.320 1196.000 374.320 ;
        RECT 4.000 336.920 1195.600 338.320 ;
        RECT 4.000 331.520 1196.000 336.920 ;
        RECT 4.400 330.120 1196.000 331.520 ;
        RECT 4.000 287.320 1196.000 330.120 ;
        RECT 4.400 285.920 1196.000 287.320 ;
        RECT 4.000 262.840 1196.000 285.920 ;
        RECT 4.000 261.440 1195.600 262.840 ;
        RECT 4.000 243.120 1196.000 261.440 ;
        RECT 4.400 241.720 1196.000 243.120 ;
        RECT 4.000 198.920 1196.000 241.720 ;
        RECT 4.400 197.520 1196.000 198.920 ;
        RECT 4.000 188.040 1196.000 197.520 ;
        RECT 4.000 186.640 1195.600 188.040 ;
        RECT 4.000 154.720 1196.000 186.640 ;
        RECT 4.400 153.320 1196.000 154.720 ;
        RECT 4.000 113.240 1196.000 153.320 ;
        RECT 4.000 111.840 1195.600 113.240 ;
        RECT 4.000 110.520 1196.000 111.840 ;
        RECT 4.400 109.120 1196.000 110.520 ;
        RECT 4.000 66.320 1196.000 109.120 ;
        RECT 4.400 64.920 1196.000 66.320 ;
        RECT 4.000 38.440 1196.000 64.920 ;
        RECT 4.000 37.040 1195.600 38.440 ;
        RECT 4.000 22.800 1196.000 37.040 ;
        RECT 4.400 21.400 1196.000 22.800 ;
        RECT 4.000 10.715 1196.000 21.400 ;
      LAYER met4 ;
        RECT 95.055 15.815 97.440 1480.185 ;
        RECT 99.840 15.815 174.240 1480.185 ;
        RECT 176.640 15.815 251.040 1480.185 ;
        RECT 253.440 15.815 327.840 1480.185 ;
        RECT 330.240 15.815 404.640 1480.185 ;
        RECT 407.040 15.815 481.440 1480.185 ;
        RECT 483.840 15.815 558.240 1480.185 ;
        RECT 560.640 15.815 635.040 1480.185 ;
        RECT 637.440 15.815 711.840 1480.185 ;
        RECT 714.240 15.815 788.640 1480.185 ;
        RECT 791.040 15.815 865.440 1480.185 ;
        RECT 867.840 15.815 942.240 1480.185 ;
        RECT 944.640 15.815 1019.040 1480.185 ;
        RECT 1021.440 15.815 1095.840 1480.185 ;
        RECT 1098.240 15.815 1172.640 1480.185 ;
        RECT 1175.040 15.815 1177.305 1480.185 ;
  END
END custom_sram
END LIBRARY

