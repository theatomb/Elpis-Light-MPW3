VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 0.000 1301.710 4.000 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.160 4.000 1349.760 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1241.040 1500.000 1241.640 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1274.360 1500.000 1274.960 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.930 0.000 1336.210 4.000 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.630 1496.000 1218.910 1500.000 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1291.360 1500.000 1291.960 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1324.680 1500.000 1325.280 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.650 1496.000 1235.930 1500.000 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 1496.000 1269.970 1500.000 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.710 1496.000 1286.990 1500.000 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 1496.000 1321.030 1500.000 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.840 4.000 1367.440 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.770 1496.000 1338.050 1500.000 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.930 0.000 1405.210 4.000 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.950 0.000 1422.230 4.000 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 4.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1407.640 1500.000 1408.240 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1419.880 4.000 1420.480 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1437.560 4.000 1438.160 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.450 0.000 1456.730 4.000 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1440.960 1500.000 1441.560 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1457.960 1500.000 1458.560 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.870 1496.000 1423.150 1500.000 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.920 4.000 1473.520 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1490.600 4.000 1491.200 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1491.280 1500.000 1491.880 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 208.120 1500.000 208.720 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 1496.000 332.490 1500.000 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 1496.000 400.570 1500.000 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 1496.000 434.610 1500.000 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 324.400 1500.000 325.000 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 357.720 1500.000 358.320 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 1496.000 536.730 1500.000 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 1496.000 553.750 1500.000 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 1496.000 587.790 1500.000 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 491.000 1500.000 491.600 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 1496.000 622.290 1500.000 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 1496.000 656.330 1500.000 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 541.320 1500.000 541.920 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 574.640 1500.000 575.240 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 4.000 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 1496.000 724.410 1500.000 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 766.400 4.000 767.000 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 590.960 1500.000 591.560 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 624.280 1500.000 624.880 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.080 4.000 784.680 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 4.000 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 641.280 1500.000 641.880 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 1496.000 758.450 1500.000 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.800 4.000 855.400 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 0.000 836.190 4.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 657.600 1500.000 658.200 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 674.600 1500.000 675.200 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 872.480 4.000 873.080 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 1496.000 809.510 1500.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 1496.000 110.770 1500.000 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 1496.000 843.550 1500.000 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 707.920 1500.000 708.520 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 741.240 1500.000 741.840 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 774.560 1500.000 775.160 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 807.880 1500.000 808.480 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 925.520 4.000 926.120 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.200 4.000 943.800 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.880 4.000 961.480 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 1496.000 894.610 1500.000 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 91.160 1500.000 91.760 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 824.880 1500.000 825.480 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 841.200 1500.000 841.800 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 874.520 1500.000 875.120 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.930 0.000 991.210 4.000 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 1496.000 929.110 1500.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 891.520 1500.000 892.120 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.430 0.000 1025.710 4.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.920 4.000 1014.520 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 907.840 1500.000 908.440 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.450 0.000 1042.730 4.000 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 1496.000 127.790 1500.000 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.930 0.000 1060.210 4.000 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 941.160 1500.000 941.760 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.280 4.000 1049.880 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 958.160 1500.000 958.760 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 991.480 1500.000 992.080 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.450 0.000 1111.730 4.000 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1024.800 1500.000 1025.400 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1041.120 1500.000 1041.720 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.000 4.000 1120.600 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.930 1496.000 1014.210 1500.000 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1058.120 1500.000 1058.720 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 1496.000 1031.230 1500.000 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 0.000 1146.230 4.000 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 1496.000 1048.250 1500.000 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 1496.000 1065.270 1500.000 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1091.440 1500.000 1092.040 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 1496.000 1099.310 1500.000 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.430 0.000 1163.710 4.000 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1260.760 4.000 1261.360 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.450 0.000 1180.730 4.000 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1296.120 4.000 1296.720 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1124.760 1500.000 1125.360 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.050 1496.000 1116.330 1500.000 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.090 1496.000 1150.370 1500.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1158.080 1500.000 1158.680 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 0.000 1249.730 4.000 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1313.800 4.000 1314.400 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.130 1496.000 1184.410 1500.000 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1174.400 1500.000 1175.000 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1331.480 4.000 1332.080 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 141.480 1500.000 142.080 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 24.520 1500.000 25.120 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 1496.000 280.970 1500.000 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 241.440 1500.000 242.040 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 274.760 1500.000 275.360 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 291.080 1500.000 291.680 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 374.720 1500.000 375.320 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 1496.000 485.670 1500.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 1496.000 570.770 1500.000 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 424.360 1500.000 424.960 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 457.680 1500.000 458.280 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 1496.000 639.310 1500.000 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 1496.000 673.350 1500.000 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1496.000 212.890 1500.000 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 157.800 1500.000 158.400 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 1496.000 42.690 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 1496.000 93.750 1500.000 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 1496.000 76.730 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 8.200 1500.000 8.800 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 1496.000 59.710 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 191.120 1500.000 191.720 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 224.440 1500.000 225.040 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 257.760 1500.000 258.360 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 1496.000 349.510 1500.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 308.080 1500.000 308.680 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 41.520 1500.000 42.120 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 108.160 1500.000 108.760 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 1496.000 161.830 1500.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 1496.000 229.910 1500.000 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.450 0.000 1318.730 4.000 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1224.720 1500.000 1225.320 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1258.040 1500.000 1258.640 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 1496.000 1201.430 1500.000 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 0.000 1370.710 4.000 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1307.680 1500.000 1308.280 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1341.000 1500.000 1341.600 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 1496.000 1252.950 1500.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1358.000 1500.000 1358.600 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.730 1496.000 1304.010 1500.000 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1374.320 1500.000 1374.920 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1391.320 1500.000 1391.920 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.450 0.000 1387.730 4.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1384.520 4.000 1385.120 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1402.200 4.000 1402.800 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.790 1496.000 1355.070 1500.000 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 1496.000 1372.090 1500.000 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1424.640 1500.000 1425.240 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.830 1496.000 1389.110 1500.000 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.850 1496.000 1406.130 1500.000 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 0.000 1474.210 4.000 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1474.280 1500.000 1474.880 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 1496.000 1440.170 1500.000 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.910 1496.000 1457.190 1500.000 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.930 1496.000 1474.210 1500.000 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 1496.000 1491.230 1500.000 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 1496.000 297.990 1500.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 1496.000 315.470 1500.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 1496.000 451.630 1500.000 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 391.040 1500.000 391.640 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 1496.000 502.690 1500.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 408.040 1500.000 408.640 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 1496.000 604.810 1500.000 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 524.320 1500.000 524.920 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 1496.000 690.370 1500.000 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 1496.000 707.390 1500.000 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 607.960 1500.000 608.560 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 0.000 767.190 4.000 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 1496.000 741.430 1500.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.760 4.000 802.360 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 57.840 1500.000 58.440 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.120 4.000 837.720 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 0.000 801.690 4.000 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 1496.000 775.470 1500.000 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 1496.000 792.490 1500.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 690.920 1500.000 691.520 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.160 4.000 890.760 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 1496.000 826.530 1500.000 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 0.000 887.710 4.000 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 724.240 1500.000 724.840 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 758.240 1500.000 758.840 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 1496.000 860.570 1500.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 791.560 1500.000 792.160 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 0.000 922.210 4.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 0.000 939.690 4.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 1496.000 877.590 1500.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 978.560 4.000 979.160 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 1496.000 912.090 1500.000 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 858.200 1500.000 858.800 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.910 0.000 974.190 4.000 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 0.000 1008.690 4.000 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.850 1496.000 946.130 1500.000 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 1496.000 963.150 1500.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1031.600 4.000 1032.200 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 924.840 1500.000 925.440 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 1496.000 980.170 1500.000 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 0.000 1077.230 4.000 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.430 0.000 1094.710 4.000 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.960 4.000 1067.560 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 974.480 1500.000 975.080 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 1496.000 997.190 1500.000 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1007.800 1500.000 1008.400 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1102.320 4.000 1102.920 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.000 4.000 1137.600 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 4.000 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 1496.000 178.850 1500.000 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1074.440 1500.000 1075.040 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.680 4.000 1155.280 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1172.360 4.000 1172.960 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.720 4.000 1208.320 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 1496.000 1082.290 1500.000 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1225.400 4.000 1226.000 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.080 4.000 1243.680 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1107.760 1500.000 1108.360 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1278.440 4.000 1279.040 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 124.480 1500.000 125.080 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 0.000 1198.210 4.000 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1141.080 1500.000 1141.680 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.070 1496.000 1133.350 1500.000 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.950 0.000 1215.230 4.000 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.430 0.000 1232.710 4.000 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.110 1496.000 1167.390 1500.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.930 0.000 1267.210 4.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.950 0.000 1284.230 4.000 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1191.400 1500.000 1192.000 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1207.720 1500.000 1208.320 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 1496.000 246.930 1500.000 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 1496.000 8.650 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 1496.000 25.670 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 174.800 1500.000 175.400 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 1496.000 366.530 1500.000 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 1496.000 383.550 1500.000 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 1496.000 417.590 1500.000 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 341.400 1500.000 342.000 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 1496.000 468.650 1500.000 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 1496.000 519.710 1500.000 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 441.360 1500.000 441.960 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 474.680 1500.000 475.280 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 508.000 1500.000 508.600 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 557.640 1500.000 558.240 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 74.840 1500.000 75.440 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 1496.000 144.810 1500.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 1496.000 195.870 1500.000 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 1496.000 263.950 1500.000 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1494.855 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.915 1489.840 ;
      LAYER met2 ;
        RECT 6.990 1495.720 8.090 1496.410 ;
        RECT 8.930 1495.720 25.110 1496.410 ;
        RECT 25.950 1495.720 42.130 1496.410 ;
        RECT 42.970 1495.720 59.150 1496.410 ;
        RECT 59.990 1495.720 76.170 1496.410 ;
        RECT 77.010 1495.720 93.190 1496.410 ;
        RECT 94.030 1495.720 110.210 1496.410 ;
        RECT 111.050 1495.720 127.230 1496.410 ;
        RECT 128.070 1495.720 144.250 1496.410 ;
        RECT 145.090 1495.720 161.270 1496.410 ;
        RECT 162.110 1495.720 178.290 1496.410 ;
        RECT 179.130 1495.720 195.310 1496.410 ;
        RECT 196.150 1495.720 212.330 1496.410 ;
        RECT 213.170 1495.720 229.350 1496.410 ;
        RECT 230.190 1495.720 246.370 1496.410 ;
        RECT 247.210 1495.720 263.390 1496.410 ;
        RECT 264.230 1495.720 280.410 1496.410 ;
        RECT 281.250 1495.720 297.430 1496.410 ;
        RECT 298.270 1495.720 314.910 1496.410 ;
        RECT 315.750 1495.720 331.930 1496.410 ;
        RECT 332.770 1495.720 348.950 1496.410 ;
        RECT 349.790 1495.720 365.970 1496.410 ;
        RECT 366.810 1495.720 382.990 1496.410 ;
        RECT 383.830 1495.720 400.010 1496.410 ;
        RECT 400.850 1495.720 417.030 1496.410 ;
        RECT 417.870 1495.720 434.050 1496.410 ;
        RECT 434.890 1495.720 451.070 1496.410 ;
        RECT 451.910 1495.720 468.090 1496.410 ;
        RECT 468.930 1495.720 485.110 1496.410 ;
        RECT 485.950 1495.720 502.130 1496.410 ;
        RECT 502.970 1495.720 519.150 1496.410 ;
        RECT 519.990 1495.720 536.170 1496.410 ;
        RECT 537.010 1495.720 553.190 1496.410 ;
        RECT 554.030 1495.720 570.210 1496.410 ;
        RECT 571.050 1495.720 587.230 1496.410 ;
        RECT 588.070 1495.720 604.250 1496.410 ;
        RECT 605.090 1495.720 621.730 1496.410 ;
        RECT 622.570 1495.720 638.750 1496.410 ;
        RECT 639.590 1495.720 655.770 1496.410 ;
        RECT 656.610 1495.720 672.790 1496.410 ;
        RECT 673.630 1495.720 689.810 1496.410 ;
        RECT 690.650 1495.720 706.830 1496.410 ;
        RECT 707.670 1495.720 723.850 1496.410 ;
        RECT 724.690 1495.720 740.870 1496.410 ;
        RECT 741.710 1495.720 757.890 1496.410 ;
        RECT 758.730 1495.720 774.910 1496.410 ;
        RECT 775.750 1495.720 791.930 1496.410 ;
        RECT 792.770 1495.720 808.950 1496.410 ;
        RECT 809.790 1495.720 825.970 1496.410 ;
        RECT 826.810 1495.720 842.990 1496.410 ;
        RECT 843.830 1495.720 860.010 1496.410 ;
        RECT 860.850 1495.720 877.030 1496.410 ;
        RECT 877.870 1495.720 894.050 1496.410 ;
        RECT 894.890 1495.720 911.530 1496.410 ;
        RECT 912.370 1495.720 928.550 1496.410 ;
        RECT 929.390 1495.720 945.570 1496.410 ;
        RECT 946.410 1495.720 962.590 1496.410 ;
        RECT 963.430 1495.720 979.610 1496.410 ;
        RECT 980.450 1495.720 996.630 1496.410 ;
        RECT 997.470 1495.720 1013.650 1496.410 ;
        RECT 1014.490 1495.720 1030.670 1496.410 ;
        RECT 1031.510 1495.720 1047.690 1496.410 ;
        RECT 1048.530 1495.720 1064.710 1496.410 ;
        RECT 1065.550 1495.720 1081.730 1496.410 ;
        RECT 1082.570 1495.720 1098.750 1496.410 ;
        RECT 1099.590 1495.720 1115.770 1496.410 ;
        RECT 1116.610 1495.720 1132.790 1496.410 ;
        RECT 1133.630 1495.720 1149.810 1496.410 ;
        RECT 1150.650 1495.720 1166.830 1496.410 ;
        RECT 1167.670 1495.720 1183.850 1496.410 ;
        RECT 1184.690 1495.720 1200.870 1496.410 ;
        RECT 1201.710 1495.720 1218.350 1496.410 ;
        RECT 1219.190 1495.720 1235.370 1496.410 ;
        RECT 1236.210 1495.720 1252.390 1496.410 ;
        RECT 1253.230 1495.720 1269.410 1496.410 ;
        RECT 1270.250 1495.720 1286.430 1496.410 ;
        RECT 1287.270 1495.720 1303.450 1496.410 ;
        RECT 1304.290 1495.720 1320.470 1496.410 ;
        RECT 1321.310 1495.720 1337.490 1496.410 ;
        RECT 1338.330 1495.720 1354.510 1496.410 ;
        RECT 1355.350 1495.720 1371.530 1496.410 ;
        RECT 1372.370 1495.720 1388.550 1496.410 ;
        RECT 1389.390 1495.720 1405.570 1496.410 ;
        RECT 1406.410 1495.720 1422.590 1496.410 ;
        RECT 1423.430 1495.720 1439.610 1496.410 ;
        RECT 1440.450 1495.720 1456.630 1496.410 ;
        RECT 1457.470 1495.720 1473.650 1496.410 ;
        RECT 1474.490 1495.720 1490.670 1496.410 ;
        RECT 6.990 4.280 1491.220 1495.720 ;
        RECT 6.990 3.670 8.090 4.280 ;
        RECT 8.930 3.670 25.110 4.280 ;
        RECT 25.950 3.670 42.130 4.280 ;
        RECT 42.970 3.670 59.610 4.280 ;
        RECT 60.450 3.670 76.630 4.280 ;
        RECT 77.470 3.670 94.110 4.280 ;
        RECT 94.950 3.670 111.130 4.280 ;
        RECT 111.970 3.670 128.610 4.280 ;
        RECT 129.450 3.670 145.630 4.280 ;
        RECT 146.470 3.670 163.110 4.280 ;
        RECT 163.950 3.670 180.130 4.280 ;
        RECT 180.970 3.670 197.610 4.280 ;
        RECT 198.450 3.670 214.630 4.280 ;
        RECT 215.470 3.670 232.110 4.280 ;
        RECT 232.950 3.670 249.130 4.280 ;
        RECT 249.970 3.670 266.610 4.280 ;
        RECT 267.450 3.670 283.630 4.280 ;
        RECT 284.470 3.670 301.110 4.280 ;
        RECT 301.950 3.670 318.130 4.280 ;
        RECT 318.970 3.670 335.610 4.280 ;
        RECT 336.450 3.670 352.630 4.280 ;
        RECT 353.470 3.670 370.110 4.280 ;
        RECT 370.950 3.670 387.130 4.280 ;
        RECT 387.970 3.670 404.610 4.280 ;
        RECT 405.450 3.670 421.630 4.280 ;
        RECT 422.470 3.670 439.110 4.280 ;
        RECT 439.950 3.670 456.130 4.280 ;
        RECT 456.970 3.670 473.610 4.280 ;
        RECT 474.450 3.670 490.630 4.280 ;
        RECT 491.470 3.670 508.110 4.280 ;
        RECT 508.950 3.670 525.130 4.280 ;
        RECT 525.970 3.670 542.150 4.280 ;
        RECT 542.990 3.670 559.630 4.280 ;
        RECT 560.470 3.670 576.650 4.280 ;
        RECT 577.490 3.670 594.130 4.280 ;
        RECT 594.970 3.670 611.150 4.280 ;
        RECT 611.990 3.670 628.630 4.280 ;
        RECT 629.470 3.670 645.650 4.280 ;
        RECT 646.490 3.670 663.130 4.280 ;
        RECT 663.970 3.670 680.150 4.280 ;
        RECT 680.990 3.670 697.630 4.280 ;
        RECT 698.470 3.670 714.650 4.280 ;
        RECT 715.490 3.670 732.130 4.280 ;
        RECT 732.970 3.670 749.150 4.280 ;
        RECT 749.990 3.670 766.630 4.280 ;
        RECT 767.470 3.670 783.650 4.280 ;
        RECT 784.490 3.670 801.130 4.280 ;
        RECT 801.970 3.670 818.150 4.280 ;
        RECT 818.990 3.670 835.630 4.280 ;
        RECT 836.470 3.670 852.650 4.280 ;
        RECT 853.490 3.670 870.130 4.280 ;
        RECT 870.970 3.670 887.150 4.280 ;
        RECT 887.990 3.670 904.630 4.280 ;
        RECT 905.470 3.670 921.650 4.280 ;
        RECT 922.490 3.670 939.130 4.280 ;
        RECT 939.970 3.670 956.150 4.280 ;
        RECT 956.990 3.670 973.630 4.280 ;
        RECT 974.470 3.670 990.650 4.280 ;
        RECT 991.490 3.670 1008.130 4.280 ;
        RECT 1008.970 3.670 1025.150 4.280 ;
        RECT 1025.990 3.670 1042.170 4.280 ;
        RECT 1043.010 3.670 1059.650 4.280 ;
        RECT 1060.490 3.670 1076.670 4.280 ;
        RECT 1077.510 3.670 1094.150 4.280 ;
        RECT 1094.990 3.670 1111.170 4.280 ;
        RECT 1112.010 3.670 1128.650 4.280 ;
        RECT 1129.490 3.670 1145.670 4.280 ;
        RECT 1146.510 3.670 1163.150 4.280 ;
        RECT 1163.990 3.670 1180.170 4.280 ;
        RECT 1181.010 3.670 1197.650 4.280 ;
        RECT 1198.490 3.670 1214.670 4.280 ;
        RECT 1215.510 3.670 1232.150 4.280 ;
        RECT 1232.990 3.670 1249.170 4.280 ;
        RECT 1250.010 3.670 1266.650 4.280 ;
        RECT 1267.490 3.670 1283.670 4.280 ;
        RECT 1284.510 3.670 1301.150 4.280 ;
        RECT 1301.990 3.670 1318.170 4.280 ;
        RECT 1319.010 3.670 1335.650 4.280 ;
        RECT 1336.490 3.670 1352.670 4.280 ;
        RECT 1353.510 3.670 1370.150 4.280 ;
        RECT 1370.990 3.670 1387.170 4.280 ;
        RECT 1388.010 3.670 1404.650 4.280 ;
        RECT 1405.490 3.670 1421.670 4.280 ;
        RECT 1422.510 3.670 1439.150 4.280 ;
        RECT 1439.990 3.670 1456.170 4.280 ;
        RECT 1457.010 3.670 1473.650 4.280 ;
        RECT 1474.490 3.670 1490.670 4.280 ;
      LAYER met3 ;
        RECT 4.000 1491.600 1495.600 1491.745 ;
        RECT 4.400 1490.880 1495.600 1491.600 ;
        RECT 4.400 1490.200 1496.000 1490.880 ;
        RECT 4.000 1475.280 1496.000 1490.200 ;
        RECT 4.000 1473.920 1495.600 1475.280 ;
        RECT 4.400 1473.880 1495.600 1473.920 ;
        RECT 4.400 1472.520 1496.000 1473.880 ;
        RECT 4.000 1458.960 1496.000 1472.520 ;
        RECT 4.000 1457.560 1495.600 1458.960 ;
        RECT 4.000 1456.240 1496.000 1457.560 ;
        RECT 4.400 1454.840 1496.000 1456.240 ;
        RECT 4.000 1441.960 1496.000 1454.840 ;
        RECT 4.000 1440.560 1495.600 1441.960 ;
        RECT 4.000 1438.560 1496.000 1440.560 ;
        RECT 4.400 1437.160 1496.000 1438.560 ;
        RECT 4.000 1425.640 1496.000 1437.160 ;
        RECT 4.000 1424.240 1495.600 1425.640 ;
        RECT 4.000 1420.880 1496.000 1424.240 ;
        RECT 4.400 1419.480 1496.000 1420.880 ;
        RECT 4.000 1408.640 1496.000 1419.480 ;
        RECT 4.000 1407.240 1495.600 1408.640 ;
        RECT 4.000 1403.200 1496.000 1407.240 ;
        RECT 4.400 1401.800 1496.000 1403.200 ;
        RECT 4.000 1392.320 1496.000 1401.800 ;
        RECT 4.000 1390.920 1495.600 1392.320 ;
        RECT 4.000 1385.520 1496.000 1390.920 ;
        RECT 4.400 1384.120 1496.000 1385.520 ;
        RECT 4.000 1375.320 1496.000 1384.120 ;
        RECT 4.000 1373.920 1495.600 1375.320 ;
        RECT 4.000 1367.840 1496.000 1373.920 ;
        RECT 4.400 1366.440 1496.000 1367.840 ;
        RECT 4.000 1359.000 1496.000 1366.440 ;
        RECT 4.000 1357.600 1495.600 1359.000 ;
        RECT 4.000 1350.160 1496.000 1357.600 ;
        RECT 4.400 1348.760 1496.000 1350.160 ;
        RECT 4.000 1342.000 1496.000 1348.760 ;
        RECT 4.000 1340.600 1495.600 1342.000 ;
        RECT 4.000 1332.480 1496.000 1340.600 ;
        RECT 4.400 1331.080 1496.000 1332.480 ;
        RECT 4.000 1325.680 1496.000 1331.080 ;
        RECT 4.000 1324.280 1495.600 1325.680 ;
        RECT 4.000 1314.800 1496.000 1324.280 ;
        RECT 4.400 1313.400 1496.000 1314.800 ;
        RECT 4.000 1308.680 1496.000 1313.400 ;
        RECT 4.000 1307.280 1495.600 1308.680 ;
        RECT 4.000 1297.120 1496.000 1307.280 ;
        RECT 4.400 1295.720 1496.000 1297.120 ;
        RECT 4.000 1292.360 1496.000 1295.720 ;
        RECT 4.000 1290.960 1495.600 1292.360 ;
        RECT 4.000 1279.440 1496.000 1290.960 ;
        RECT 4.400 1278.040 1496.000 1279.440 ;
        RECT 4.000 1275.360 1496.000 1278.040 ;
        RECT 4.000 1273.960 1495.600 1275.360 ;
        RECT 4.000 1261.760 1496.000 1273.960 ;
        RECT 4.400 1260.360 1496.000 1261.760 ;
        RECT 4.000 1259.040 1496.000 1260.360 ;
        RECT 4.000 1257.640 1495.600 1259.040 ;
        RECT 4.000 1244.080 1496.000 1257.640 ;
        RECT 4.400 1242.680 1496.000 1244.080 ;
        RECT 4.000 1242.040 1496.000 1242.680 ;
        RECT 4.000 1240.640 1495.600 1242.040 ;
        RECT 4.000 1226.400 1496.000 1240.640 ;
        RECT 4.400 1225.720 1496.000 1226.400 ;
        RECT 4.400 1225.000 1495.600 1225.720 ;
        RECT 4.000 1224.320 1495.600 1225.000 ;
        RECT 4.000 1208.720 1496.000 1224.320 ;
        RECT 4.400 1207.320 1495.600 1208.720 ;
        RECT 4.000 1192.400 1496.000 1207.320 ;
        RECT 4.000 1191.040 1495.600 1192.400 ;
        RECT 4.400 1191.000 1495.600 1191.040 ;
        RECT 4.400 1189.640 1496.000 1191.000 ;
        RECT 4.000 1175.400 1496.000 1189.640 ;
        RECT 4.000 1174.000 1495.600 1175.400 ;
        RECT 4.000 1173.360 1496.000 1174.000 ;
        RECT 4.400 1171.960 1496.000 1173.360 ;
        RECT 4.000 1159.080 1496.000 1171.960 ;
        RECT 4.000 1157.680 1495.600 1159.080 ;
        RECT 4.000 1155.680 1496.000 1157.680 ;
        RECT 4.400 1154.280 1496.000 1155.680 ;
        RECT 4.000 1142.080 1496.000 1154.280 ;
        RECT 4.000 1140.680 1495.600 1142.080 ;
        RECT 4.000 1138.000 1496.000 1140.680 ;
        RECT 4.400 1136.600 1496.000 1138.000 ;
        RECT 4.000 1125.760 1496.000 1136.600 ;
        RECT 4.000 1124.360 1495.600 1125.760 ;
        RECT 4.000 1121.000 1496.000 1124.360 ;
        RECT 4.400 1119.600 1496.000 1121.000 ;
        RECT 4.000 1108.760 1496.000 1119.600 ;
        RECT 4.000 1107.360 1495.600 1108.760 ;
        RECT 4.000 1103.320 1496.000 1107.360 ;
        RECT 4.400 1101.920 1496.000 1103.320 ;
        RECT 4.000 1092.440 1496.000 1101.920 ;
        RECT 4.000 1091.040 1495.600 1092.440 ;
        RECT 4.000 1085.640 1496.000 1091.040 ;
        RECT 4.400 1084.240 1496.000 1085.640 ;
        RECT 4.000 1075.440 1496.000 1084.240 ;
        RECT 4.000 1074.040 1495.600 1075.440 ;
        RECT 4.000 1067.960 1496.000 1074.040 ;
        RECT 4.400 1066.560 1496.000 1067.960 ;
        RECT 4.000 1059.120 1496.000 1066.560 ;
        RECT 4.000 1057.720 1495.600 1059.120 ;
        RECT 4.000 1050.280 1496.000 1057.720 ;
        RECT 4.400 1048.880 1496.000 1050.280 ;
        RECT 4.000 1042.120 1496.000 1048.880 ;
        RECT 4.000 1040.720 1495.600 1042.120 ;
        RECT 4.000 1032.600 1496.000 1040.720 ;
        RECT 4.400 1031.200 1496.000 1032.600 ;
        RECT 4.000 1025.800 1496.000 1031.200 ;
        RECT 4.000 1024.400 1495.600 1025.800 ;
        RECT 4.000 1014.920 1496.000 1024.400 ;
        RECT 4.400 1013.520 1496.000 1014.920 ;
        RECT 4.000 1008.800 1496.000 1013.520 ;
        RECT 4.000 1007.400 1495.600 1008.800 ;
        RECT 4.000 997.240 1496.000 1007.400 ;
        RECT 4.400 995.840 1496.000 997.240 ;
        RECT 4.000 992.480 1496.000 995.840 ;
        RECT 4.000 991.080 1495.600 992.480 ;
        RECT 4.000 979.560 1496.000 991.080 ;
        RECT 4.400 978.160 1496.000 979.560 ;
        RECT 4.000 975.480 1496.000 978.160 ;
        RECT 4.000 974.080 1495.600 975.480 ;
        RECT 4.000 961.880 1496.000 974.080 ;
        RECT 4.400 960.480 1496.000 961.880 ;
        RECT 4.000 959.160 1496.000 960.480 ;
        RECT 4.000 957.760 1495.600 959.160 ;
        RECT 4.000 944.200 1496.000 957.760 ;
        RECT 4.400 942.800 1496.000 944.200 ;
        RECT 4.000 942.160 1496.000 942.800 ;
        RECT 4.000 940.760 1495.600 942.160 ;
        RECT 4.000 926.520 1496.000 940.760 ;
        RECT 4.400 925.840 1496.000 926.520 ;
        RECT 4.400 925.120 1495.600 925.840 ;
        RECT 4.000 924.440 1495.600 925.120 ;
        RECT 4.000 908.840 1496.000 924.440 ;
        RECT 4.400 907.440 1495.600 908.840 ;
        RECT 4.000 892.520 1496.000 907.440 ;
        RECT 4.000 891.160 1495.600 892.520 ;
        RECT 4.400 891.120 1495.600 891.160 ;
        RECT 4.400 889.760 1496.000 891.120 ;
        RECT 4.000 875.520 1496.000 889.760 ;
        RECT 4.000 874.120 1495.600 875.520 ;
        RECT 4.000 873.480 1496.000 874.120 ;
        RECT 4.400 872.080 1496.000 873.480 ;
        RECT 4.000 859.200 1496.000 872.080 ;
        RECT 4.000 857.800 1495.600 859.200 ;
        RECT 4.000 855.800 1496.000 857.800 ;
        RECT 4.400 854.400 1496.000 855.800 ;
        RECT 4.000 842.200 1496.000 854.400 ;
        RECT 4.000 840.800 1495.600 842.200 ;
        RECT 4.000 838.120 1496.000 840.800 ;
        RECT 4.400 836.720 1496.000 838.120 ;
        RECT 4.000 825.880 1496.000 836.720 ;
        RECT 4.000 824.480 1495.600 825.880 ;
        RECT 4.000 820.440 1496.000 824.480 ;
        RECT 4.400 819.040 1496.000 820.440 ;
        RECT 4.000 808.880 1496.000 819.040 ;
        RECT 4.000 807.480 1495.600 808.880 ;
        RECT 4.000 802.760 1496.000 807.480 ;
        RECT 4.400 801.360 1496.000 802.760 ;
        RECT 4.000 792.560 1496.000 801.360 ;
        RECT 4.000 791.160 1495.600 792.560 ;
        RECT 4.000 785.080 1496.000 791.160 ;
        RECT 4.400 783.680 1496.000 785.080 ;
        RECT 4.000 775.560 1496.000 783.680 ;
        RECT 4.000 774.160 1495.600 775.560 ;
        RECT 4.000 767.400 1496.000 774.160 ;
        RECT 4.400 766.000 1496.000 767.400 ;
        RECT 4.000 759.240 1496.000 766.000 ;
        RECT 4.000 757.840 1495.600 759.240 ;
        RECT 4.000 750.400 1496.000 757.840 ;
        RECT 4.400 749.000 1496.000 750.400 ;
        RECT 4.000 742.240 1496.000 749.000 ;
        RECT 4.000 740.840 1495.600 742.240 ;
        RECT 4.000 732.720 1496.000 740.840 ;
        RECT 4.400 731.320 1496.000 732.720 ;
        RECT 4.000 725.240 1496.000 731.320 ;
        RECT 4.000 723.840 1495.600 725.240 ;
        RECT 4.000 715.040 1496.000 723.840 ;
        RECT 4.400 713.640 1496.000 715.040 ;
        RECT 4.000 708.920 1496.000 713.640 ;
        RECT 4.000 707.520 1495.600 708.920 ;
        RECT 4.000 697.360 1496.000 707.520 ;
        RECT 4.400 695.960 1496.000 697.360 ;
        RECT 4.000 691.920 1496.000 695.960 ;
        RECT 4.000 690.520 1495.600 691.920 ;
        RECT 4.000 679.680 1496.000 690.520 ;
        RECT 4.400 678.280 1496.000 679.680 ;
        RECT 4.000 675.600 1496.000 678.280 ;
        RECT 4.000 674.200 1495.600 675.600 ;
        RECT 4.000 662.000 1496.000 674.200 ;
        RECT 4.400 660.600 1496.000 662.000 ;
        RECT 4.000 658.600 1496.000 660.600 ;
        RECT 4.000 657.200 1495.600 658.600 ;
        RECT 4.000 644.320 1496.000 657.200 ;
        RECT 4.400 642.920 1496.000 644.320 ;
        RECT 4.000 642.280 1496.000 642.920 ;
        RECT 4.000 640.880 1495.600 642.280 ;
        RECT 4.000 626.640 1496.000 640.880 ;
        RECT 4.400 625.280 1496.000 626.640 ;
        RECT 4.400 625.240 1495.600 625.280 ;
        RECT 4.000 623.880 1495.600 625.240 ;
        RECT 4.000 608.960 1496.000 623.880 ;
        RECT 4.400 607.560 1495.600 608.960 ;
        RECT 4.000 591.960 1496.000 607.560 ;
        RECT 4.000 591.280 1495.600 591.960 ;
        RECT 4.400 590.560 1495.600 591.280 ;
        RECT 4.400 589.880 1496.000 590.560 ;
        RECT 4.000 575.640 1496.000 589.880 ;
        RECT 4.000 574.240 1495.600 575.640 ;
        RECT 4.000 573.600 1496.000 574.240 ;
        RECT 4.400 572.200 1496.000 573.600 ;
        RECT 4.000 558.640 1496.000 572.200 ;
        RECT 4.000 557.240 1495.600 558.640 ;
        RECT 4.000 555.920 1496.000 557.240 ;
        RECT 4.400 554.520 1496.000 555.920 ;
        RECT 4.000 542.320 1496.000 554.520 ;
        RECT 4.000 540.920 1495.600 542.320 ;
        RECT 4.000 538.240 1496.000 540.920 ;
        RECT 4.400 536.840 1496.000 538.240 ;
        RECT 4.000 525.320 1496.000 536.840 ;
        RECT 4.000 523.920 1495.600 525.320 ;
        RECT 4.000 520.560 1496.000 523.920 ;
        RECT 4.400 519.160 1496.000 520.560 ;
        RECT 4.000 509.000 1496.000 519.160 ;
        RECT 4.000 507.600 1495.600 509.000 ;
        RECT 4.000 502.880 1496.000 507.600 ;
        RECT 4.400 501.480 1496.000 502.880 ;
        RECT 4.000 492.000 1496.000 501.480 ;
        RECT 4.000 490.600 1495.600 492.000 ;
        RECT 4.000 485.200 1496.000 490.600 ;
        RECT 4.400 483.800 1496.000 485.200 ;
        RECT 4.000 475.680 1496.000 483.800 ;
        RECT 4.000 474.280 1495.600 475.680 ;
        RECT 4.000 467.520 1496.000 474.280 ;
        RECT 4.400 466.120 1496.000 467.520 ;
        RECT 4.000 458.680 1496.000 466.120 ;
        RECT 4.000 457.280 1495.600 458.680 ;
        RECT 4.000 449.840 1496.000 457.280 ;
        RECT 4.400 448.440 1496.000 449.840 ;
        RECT 4.000 442.360 1496.000 448.440 ;
        RECT 4.000 440.960 1495.600 442.360 ;
        RECT 4.000 432.160 1496.000 440.960 ;
        RECT 4.400 430.760 1496.000 432.160 ;
        RECT 4.000 425.360 1496.000 430.760 ;
        RECT 4.000 423.960 1495.600 425.360 ;
        RECT 4.000 414.480 1496.000 423.960 ;
        RECT 4.400 413.080 1496.000 414.480 ;
        RECT 4.000 409.040 1496.000 413.080 ;
        RECT 4.000 407.640 1495.600 409.040 ;
        RECT 4.000 396.800 1496.000 407.640 ;
        RECT 4.400 395.400 1496.000 396.800 ;
        RECT 4.000 392.040 1496.000 395.400 ;
        RECT 4.000 390.640 1495.600 392.040 ;
        RECT 4.000 379.800 1496.000 390.640 ;
        RECT 4.400 378.400 1496.000 379.800 ;
        RECT 4.000 375.720 1496.000 378.400 ;
        RECT 4.000 374.320 1495.600 375.720 ;
        RECT 4.000 362.120 1496.000 374.320 ;
        RECT 4.400 360.720 1496.000 362.120 ;
        RECT 4.000 358.720 1496.000 360.720 ;
        RECT 4.000 357.320 1495.600 358.720 ;
        RECT 4.000 344.440 1496.000 357.320 ;
        RECT 4.400 343.040 1496.000 344.440 ;
        RECT 4.000 342.400 1496.000 343.040 ;
        RECT 4.000 341.000 1495.600 342.400 ;
        RECT 4.000 326.760 1496.000 341.000 ;
        RECT 4.400 325.400 1496.000 326.760 ;
        RECT 4.400 325.360 1495.600 325.400 ;
        RECT 4.000 324.000 1495.600 325.360 ;
        RECT 4.000 309.080 1496.000 324.000 ;
        RECT 4.400 307.680 1495.600 309.080 ;
        RECT 4.000 292.080 1496.000 307.680 ;
        RECT 4.000 291.400 1495.600 292.080 ;
        RECT 4.400 290.680 1495.600 291.400 ;
        RECT 4.400 290.000 1496.000 290.680 ;
        RECT 4.000 275.760 1496.000 290.000 ;
        RECT 4.000 274.360 1495.600 275.760 ;
        RECT 4.000 273.720 1496.000 274.360 ;
        RECT 4.400 272.320 1496.000 273.720 ;
        RECT 4.000 258.760 1496.000 272.320 ;
        RECT 4.000 257.360 1495.600 258.760 ;
        RECT 4.000 256.040 1496.000 257.360 ;
        RECT 4.400 254.640 1496.000 256.040 ;
        RECT 4.000 242.440 1496.000 254.640 ;
        RECT 4.000 241.040 1495.600 242.440 ;
        RECT 4.000 238.360 1496.000 241.040 ;
        RECT 4.400 236.960 1496.000 238.360 ;
        RECT 4.000 225.440 1496.000 236.960 ;
        RECT 4.000 224.040 1495.600 225.440 ;
        RECT 4.000 220.680 1496.000 224.040 ;
        RECT 4.400 219.280 1496.000 220.680 ;
        RECT 4.000 209.120 1496.000 219.280 ;
        RECT 4.000 207.720 1495.600 209.120 ;
        RECT 4.000 203.000 1496.000 207.720 ;
        RECT 4.400 201.600 1496.000 203.000 ;
        RECT 4.000 192.120 1496.000 201.600 ;
        RECT 4.000 190.720 1495.600 192.120 ;
        RECT 4.000 185.320 1496.000 190.720 ;
        RECT 4.400 183.920 1496.000 185.320 ;
        RECT 4.000 175.800 1496.000 183.920 ;
        RECT 4.000 174.400 1495.600 175.800 ;
        RECT 4.000 167.640 1496.000 174.400 ;
        RECT 4.400 166.240 1496.000 167.640 ;
        RECT 4.000 158.800 1496.000 166.240 ;
        RECT 4.000 157.400 1495.600 158.800 ;
        RECT 4.000 149.960 1496.000 157.400 ;
        RECT 4.400 148.560 1496.000 149.960 ;
        RECT 4.000 142.480 1496.000 148.560 ;
        RECT 4.000 141.080 1495.600 142.480 ;
        RECT 4.000 132.280 1496.000 141.080 ;
        RECT 4.400 130.880 1496.000 132.280 ;
        RECT 4.000 125.480 1496.000 130.880 ;
        RECT 4.000 124.080 1495.600 125.480 ;
        RECT 4.000 114.600 1496.000 124.080 ;
        RECT 4.400 113.200 1496.000 114.600 ;
        RECT 4.000 109.160 1496.000 113.200 ;
        RECT 4.000 107.760 1495.600 109.160 ;
        RECT 4.000 96.920 1496.000 107.760 ;
        RECT 4.400 95.520 1496.000 96.920 ;
        RECT 4.000 92.160 1496.000 95.520 ;
        RECT 4.000 90.760 1495.600 92.160 ;
        RECT 4.000 79.240 1496.000 90.760 ;
        RECT 4.400 77.840 1496.000 79.240 ;
        RECT 4.000 75.840 1496.000 77.840 ;
        RECT 4.000 74.440 1495.600 75.840 ;
        RECT 4.000 61.560 1496.000 74.440 ;
        RECT 4.400 60.160 1496.000 61.560 ;
        RECT 4.000 58.840 1496.000 60.160 ;
        RECT 4.000 57.440 1495.600 58.840 ;
        RECT 4.000 43.880 1496.000 57.440 ;
        RECT 4.400 42.520 1496.000 43.880 ;
        RECT 4.400 42.480 1495.600 42.520 ;
        RECT 4.000 41.120 1495.600 42.480 ;
        RECT 4.000 26.200 1496.000 41.120 ;
        RECT 4.400 25.520 1496.000 26.200 ;
        RECT 4.400 24.800 1495.600 25.520 ;
        RECT 4.000 24.120 1495.600 24.800 ;
        RECT 4.000 9.200 1496.000 24.120 ;
        RECT 4.400 8.335 1495.600 9.200 ;
      LAYER met4 ;
        RECT 193.495 10.240 251.040 1480.185 ;
        RECT 253.440 10.240 327.840 1480.185 ;
        RECT 330.240 10.240 404.640 1480.185 ;
        RECT 407.040 10.240 481.440 1480.185 ;
        RECT 483.840 10.240 558.240 1480.185 ;
        RECT 560.640 10.240 635.040 1480.185 ;
        RECT 637.440 10.240 711.840 1480.185 ;
        RECT 714.240 10.240 788.640 1480.185 ;
        RECT 791.040 10.240 865.440 1480.185 ;
        RECT 867.840 10.240 942.240 1480.185 ;
        RECT 944.640 10.240 1019.040 1480.185 ;
        RECT 1021.440 10.240 1061.385 1480.185 ;
        RECT 193.495 9.695 1061.385 10.240 ;
  END
END core
END LIBRARY

