VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO custom_sram
  CLASS BLOCK ;
  FOREIGN custom_sram ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1500.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 1496.000 566.630 1500.000 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 608.640 1200.000 609.240 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.000 4.000 916.600 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 796.320 1200.000 796.920 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 983.320 1200.000 983.920 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 139.440 1200.000 140.040 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 1496.000 33.490 1500.000 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 327.120 1200.000 327.720 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 1496.000 366.530 1500.000 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END a[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END clk
  PIN csb0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END csb0_to_sram
  PIN d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END d[0]
  PIN d[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 1496.000 499.930 1500.000 ;
    END
  END d[10]
  PIN d[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 1496.000 633.330 1500.000 ;
    END
  END d[11]
  PIN d[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.800 4.000 583.400 ;
    END
  END d[12]
  PIN d[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 702.480 1200.000 703.080 ;
    END
  END d[13]
  PIN d[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END d[14]
  PIN d[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END d[15]
  PIN d[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END d[16]
  PIN d[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 889.480 1200.000 890.080 ;
    END
  END d[17]
  PIN d[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 1496.000 766.730 1500.000 ;
    END
  END d[18]
  PIN d[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 1496.000 833.430 1500.000 ;
    END
  END d[19]
  PIN d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 233.280 1200.000 233.880 ;
    END
  END d[1]
  PIN d[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 0.000 911.170 4.000 ;
    END
  END d[20]
  PIN d[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 4.000 ;
    END
  END d[21]
  PIN d[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1496.000 900.130 1500.000 ;
    END
  END d[22]
  PIN d[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 0.000 1044.570 4.000 ;
    END
  END d[23]
  PIN d[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1171.000 1200.000 1171.600 ;
    END
  END d[24]
  PIN d[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1249.200 4.000 1249.800 ;
    END
  END d[25]
  PIN d[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 0.000 1089.190 4.000 ;
    END
  END d[26]
  PIN d[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1358.680 1200.000 1359.280 ;
    END
  END d[27]
  PIN d[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.070 0.000 1133.350 4.000 ;
    END
  END d[28]
  PIN d[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 1496.000 1100.230 1500.000 ;
    END
  END d[29]
  PIN d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END d[2]
  PIN d[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END d[30]
  PIN d[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1415.800 4.000 1416.400 ;
    END
  END d[31]
  PIN d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END d[3]
  PIN d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 1496.000 166.430 1500.000 ;
    END
  END d[4]
  PIN d[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 514.800 1200.000 515.400 ;
    END
  END d[5]
  PIN d[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END d[6]
  PIN d[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 1496.000 433.230 1500.000 ;
    END
  END d[7]
  PIN d[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END d[8]
  PIN d[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END d[9]
  PIN q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 46.280 1200.000 46.880 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 1496.000 700.030 1500.000 ;
    END
  END q[11]
  PIN q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END q[12]
  PIN q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END q[13]
  PIN q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 804.480 4.000 805.080 ;
    END
  END q[14]
  PIN q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END q[15]
  PIN q[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END q[16]
  PIN q[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END q[17]
  PIN q[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1026.840 4.000 1027.440 ;
    END
  END q[18]
  PIN q[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1077.160 1200.000 1077.760 ;
    END
  END q[19]
  PIN q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END q[1]
  PIN q[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.510 0.000 955.790 4.000 ;
    END
  END q[20]
  PIN q[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1082.600 4.000 1083.200 ;
    END
  END q[21]
  PIN q[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1138.360 4.000 1138.960 ;
    END
  END q[22]
  PIN q[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END q[23]
  PIN q[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1264.840 1200.000 1265.440 ;
    END
  END q[24]
  PIN q[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 1496.000 966.830 1500.000 ;
    END
  END q[25]
  PIN q[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 1496.000 1033.530 1500.000 ;
    END
  END q[26]
  PIN q[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1304.960 4.000 1305.560 ;
    END
  END q[27]
  PIN q[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1452.520 1200.000 1453.120 ;
    END
  END q[28]
  PIN q[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.690 0.000 1177.970 4.000 ;
    END
  END q[29]
  PIN q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 1496.000 99.730 1500.000 ;
    END
  END q[2]
  PIN q[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.650 1496.000 1166.930 1500.000 ;
    END
  END q[30]
  PIN q[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1471.560 4.000 1472.160 ;
    END
  END q[31]
  PIN q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 420.960 1200.000 421.560 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 1496.000 233.130 1500.000 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1496.000 299.830 1500.000 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END q[9]
  PIN spare_wen0_to_sram
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
  END vssd1
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END we
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1196.775 1487.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 1196.835 1488.080 ;
      LAYER met2 ;
        RECT 6.990 1495.720 32.930 1496.410 ;
        RECT 33.770 1495.720 99.170 1496.410 ;
        RECT 100.010 1495.720 165.870 1496.410 ;
        RECT 166.710 1495.720 232.570 1496.410 ;
        RECT 233.410 1495.720 299.270 1496.410 ;
        RECT 300.110 1495.720 365.970 1496.410 ;
        RECT 366.810 1495.720 432.670 1496.410 ;
        RECT 433.510 1495.720 499.370 1496.410 ;
        RECT 500.210 1495.720 566.070 1496.410 ;
        RECT 566.910 1495.720 632.770 1496.410 ;
        RECT 633.610 1495.720 699.470 1496.410 ;
        RECT 700.310 1495.720 766.170 1496.410 ;
        RECT 767.010 1495.720 832.870 1496.410 ;
        RECT 833.710 1495.720 899.570 1496.410 ;
        RECT 900.410 1495.720 966.270 1496.410 ;
        RECT 967.110 1495.720 1032.970 1496.410 ;
        RECT 1033.810 1495.720 1099.670 1496.410 ;
        RECT 1100.510 1495.720 1166.370 1496.410 ;
        RECT 1167.210 1495.720 1194.990 1496.410 ;
        RECT 6.990 4.280 1194.990 1495.720 ;
        RECT 6.990 3.670 21.890 4.280 ;
        RECT 22.730 3.670 66.050 4.280 ;
        RECT 66.890 3.670 110.670 4.280 ;
        RECT 111.510 3.670 154.830 4.280 ;
        RECT 155.670 3.670 199.450 4.280 ;
        RECT 200.290 3.670 244.070 4.280 ;
        RECT 244.910 3.670 288.230 4.280 ;
        RECT 289.070 3.670 332.850 4.280 ;
        RECT 333.690 3.670 377.470 4.280 ;
        RECT 378.310 3.670 421.630 4.280 ;
        RECT 422.470 3.670 466.250 4.280 ;
        RECT 467.090 3.670 510.410 4.280 ;
        RECT 511.250 3.670 555.030 4.280 ;
        RECT 555.870 3.670 599.650 4.280 ;
        RECT 600.490 3.670 643.810 4.280 ;
        RECT 644.650 3.670 688.430 4.280 ;
        RECT 689.270 3.670 733.050 4.280 ;
        RECT 733.890 3.670 777.210 4.280 ;
        RECT 778.050 3.670 821.830 4.280 ;
        RECT 822.670 3.670 865.990 4.280 ;
        RECT 866.830 3.670 910.610 4.280 ;
        RECT 911.450 3.670 955.230 4.280 ;
        RECT 956.070 3.670 999.390 4.280 ;
        RECT 1000.230 3.670 1044.010 4.280 ;
        RECT 1044.850 3.670 1088.630 4.280 ;
        RECT 1089.470 3.670 1132.790 4.280 ;
        RECT 1133.630 3.670 1177.410 4.280 ;
        RECT 1178.250 3.670 1194.990 4.280 ;
      LAYER met3 ;
        RECT 4.000 1472.560 1196.000 1488.005 ;
        RECT 4.400 1471.160 1196.000 1472.560 ;
        RECT 4.000 1453.520 1196.000 1471.160 ;
        RECT 4.000 1452.120 1195.600 1453.520 ;
        RECT 4.000 1416.800 1196.000 1452.120 ;
        RECT 4.400 1415.400 1196.000 1416.800 ;
        RECT 4.000 1361.040 1196.000 1415.400 ;
        RECT 4.400 1359.680 1196.000 1361.040 ;
        RECT 4.400 1359.640 1195.600 1359.680 ;
        RECT 4.000 1358.280 1195.600 1359.640 ;
        RECT 4.000 1305.960 1196.000 1358.280 ;
        RECT 4.400 1304.560 1196.000 1305.960 ;
        RECT 4.000 1265.840 1196.000 1304.560 ;
        RECT 4.000 1264.440 1195.600 1265.840 ;
        RECT 4.000 1250.200 1196.000 1264.440 ;
        RECT 4.400 1248.800 1196.000 1250.200 ;
        RECT 4.000 1194.440 1196.000 1248.800 ;
        RECT 4.400 1193.040 1196.000 1194.440 ;
        RECT 4.000 1172.000 1196.000 1193.040 ;
        RECT 4.000 1170.600 1195.600 1172.000 ;
        RECT 4.000 1139.360 1196.000 1170.600 ;
        RECT 4.400 1137.960 1196.000 1139.360 ;
        RECT 4.000 1083.600 1196.000 1137.960 ;
        RECT 4.400 1082.200 1196.000 1083.600 ;
        RECT 4.000 1078.160 1196.000 1082.200 ;
        RECT 4.000 1076.760 1195.600 1078.160 ;
        RECT 4.000 1027.840 1196.000 1076.760 ;
        RECT 4.400 1026.440 1196.000 1027.840 ;
        RECT 4.000 984.320 1196.000 1026.440 ;
        RECT 4.000 982.920 1195.600 984.320 ;
        RECT 4.000 972.080 1196.000 982.920 ;
        RECT 4.400 970.680 1196.000 972.080 ;
        RECT 4.000 917.000 1196.000 970.680 ;
        RECT 4.400 915.600 1196.000 917.000 ;
        RECT 4.000 890.480 1196.000 915.600 ;
        RECT 4.000 889.080 1195.600 890.480 ;
        RECT 4.000 861.240 1196.000 889.080 ;
        RECT 4.400 859.840 1196.000 861.240 ;
        RECT 4.000 805.480 1196.000 859.840 ;
        RECT 4.400 804.080 1196.000 805.480 ;
        RECT 4.000 797.320 1196.000 804.080 ;
        RECT 4.000 795.920 1195.600 797.320 ;
        RECT 4.000 750.400 1196.000 795.920 ;
        RECT 4.400 749.000 1196.000 750.400 ;
        RECT 4.000 703.480 1196.000 749.000 ;
        RECT 4.000 702.080 1195.600 703.480 ;
        RECT 4.000 694.640 1196.000 702.080 ;
        RECT 4.400 693.240 1196.000 694.640 ;
        RECT 4.000 638.880 1196.000 693.240 ;
        RECT 4.400 637.480 1196.000 638.880 ;
        RECT 4.000 609.640 1196.000 637.480 ;
        RECT 4.000 608.240 1195.600 609.640 ;
        RECT 4.000 583.800 1196.000 608.240 ;
        RECT 4.400 582.400 1196.000 583.800 ;
        RECT 4.000 528.040 1196.000 582.400 ;
        RECT 4.400 526.640 1196.000 528.040 ;
        RECT 4.000 515.800 1196.000 526.640 ;
        RECT 4.000 514.400 1195.600 515.800 ;
        RECT 4.000 472.280 1196.000 514.400 ;
        RECT 4.400 470.880 1196.000 472.280 ;
        RECT 4.000 421.960 1196.000 470.880 ;
        RECT 4.000 420.560 1195.600 421.960 ;
        RECT 4.000 416.520 1196.000 420.560 ;
        RECT 4.400 415.120 1196.000 416.520 ;
        RECT 4.000 361.440 1196.000 415.120 ;
        RECT 4.400 360.040 1196.000 361.440 ;
        RECT 4.000 328.120 1196.000 360.040 ;
        RECT 4.000 326.720 1195.600 328.120 ;
        RECT 4.000 305.680 1196.000 326.720 ;
        RECT 4.400 304.280 1196.000 305.680 ;
        RECT 4.000 249.920 1196.000 304.280 ;
        RECT 4.400 248.520 1196.000 249.920 ;
        RECT 4.000 234.280 1196.000 248.520 ;
        RECT 4.000 232.880 1195.600 234.280 ;
        RECT 4.000 194.840 1196.000 232.880 ;
        RECT 4.400 193.440 1196.000 194.840 ;
        RECT 4.000 140.440 1196.000 193.440 ;
        RECT 4.000 139.080 1195.600 140.440 ;
        RECT 4.400 139.040 1195.600 139.080 ;
        RECT 4.400 137.680 1196.000 139.040 ;
        RECT 4.000 83.320 1196.000 137.680 ;
        RECT 4.400 81.920 1196.000 83.320 ;
        RECT 4.000 47.280 1196.000 81.920 ;
        RECT 4.000 45.880 1195.600 47.280 ;
        RECT 4.000 28.240 1196.000 45.880 ;
        RECT 4.400 26.840 1196.000 28.240 ;
        RECT 4.000 10.715 1196.000 26.840 ;
      LAYER met4 ;
        RECT 91.375 18.535 97.440 1442.785 ;
        RECT 99.840 18.535 174.240 1442.785 ;
        RECT 176.640 18.535 251.040 1442.785 ;
        RECT 253.440 18.535 327.840 1442.785 ;
        RECT 330.240 18.535 404.640 1442.785 ;
        RECT 407.040 18.535 481.440 1442.785 ;
        RECT 483.840 18.535 558.240 1442.785 ;
        RECT 560.640 18.535 635.040 1442.785 ;
        RECT 637.440 18.535 711.840 1442.785 ;
        RECT 714.240 18.535 788.640 1442.785 ;
        RECT 791.040 18.535 865.440 1442.785 ;
        RECT 867.840 18.535 942.240 1442.785 ;
        RECT 944.640 18.535 1019.040 1442.785 ;
        RECT 1021.440 18.535 1095.840 1442.785 ;
        RECT 1098.240 18.535 1172.640 1442.785 ;
        RECT 1175.040 18.535 1175.465 1442.785 ;
  END
END custom_sram
END LIBRARY

