VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 1496.000 9.570 1500.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.950 1496.000 1284.230 1500.000 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.080 4.000 1243.680 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.170 0.000 1310.450 4.000 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 4.000 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1263.480 1500.000 1264.080 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1281.160 1500.000 1281.760 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.530 1496.000 1340.810 1500.000 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.530 0.000 1340.810 4.000 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.710 0.000 1355.990 4.000 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1296.120 4.000 1296.720 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1315.840 1500.000 1316.440 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.070 0.000 1386.350 4.000 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1368.200 1500.000 1368.800 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.650 1496.000 1396.930 1500.000 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.910 1496.000 1434.190 1500.000 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.770 1496.000 1453.050 1500.000 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 1496.000 1490.770 1500.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1385.880 1500.000 1386.480 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1403.560 1500.000 1404.160 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.430 0.000 1416.710 4.000 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 199.960 1500.000 200.560 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.610 0.000 1431.890 4.000 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1384.520 4.000 1385.120 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1419.880 4.000 1420.480 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1438.240 1500.000 1438.840 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.330 0.000 1492.610 4.000 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1472.920 1500.000 1473.520 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 4.000 1455.840 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.920 4.000 1473.520 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 1496.000 346.750 1500.000 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 1496.000 421.730 1500.000 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 1496.000 140.670 1500.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 1496.000 515.570 1500.000 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 391.720 1500.000 392.320 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 1496.000 590.550 1500.000 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 444.080 1500.000 444.680 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 1496.000 665.530 1500.000 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 1496.000 159.530 1500.000 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 1496.000 703.250 1500.000 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.080 4.000 784.680 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 601.160 1500.000 601.760 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 618.160 1500.000 618.760 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 1496.000 759.370 1500.000 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 0.000 719.810 4.000 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 4.000 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 670.520 1500.000 671.120 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 1496.000 778.230 1500.000 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 0.000 795.250 4.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 688.200 1500.000 688.800 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 705.880 1500.000 706.480 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 1496.000 815.490 1500.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 77.560 1500.000 78.160 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 0.000 886.330 4.000 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 1496.000 834.350 1500.000 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 4.000 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 1496.000 853.210 1500.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 1496.000 872.070 1500.000 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 0.000 962.230 4.000 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 758.240 1500.000 758.840 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 0.000 1007.770 4.000 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 792.920 1500.000 793.520 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 925.520 4.000 926.120 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 1496.000 909.330 1500.000 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 1496.000 947.050 1500.000 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.570 0.000 1052.850 4.000 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 0.000 1068.030 4.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.880 4.000 961.480 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 0.000 1083.210 4.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 845.280 1500.000 845.880 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 0.000 1113.570 4.000 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 1496.000 215.650 1500.000 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.920 4.000 1014.520 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 1496.000 1003.170 1500.000 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1031.600 4.000 1032.200 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 1496.000 1040.430 1500.000 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.830 0.000 1159.110 4.000 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 1496.000 1059.290 1500.000 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 914.640 1500.000 915.240 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1102.320 4.000 1102.920 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.190 0.000 1189.470 4.000 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.000 4.000 1137.600 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 1496.000 1115.410 1500.000 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 984.680 1500.000 985.280 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.990 1496.000 1134.270 1500.000 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.680 4.000 1155.280 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1002.360 1500.000 1002.960 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.850 1496.000 1153.130 1500.000 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1037.040 1500.000 1037.640 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.710 1496.000 1171.990 1500.000 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1089.400 1500.000 1090.000 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1124.080 1500.000 1124.680 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.630 0.000 1264.910 4.000 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.970 1496.000 1209.250 1500.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1172.360 4.000 1172.960 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1176.440 1500.000 1177.040 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1194.120 1500.000 1194.720 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 1496.000 1246.970 1500.000 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.040 4.000 1190.640 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1228.800 1500.000 1229.400 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 1496.000 271.770 1500.000 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 216.960 1500.000 217.560 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 1496.000 403.330 1500.000 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 1496.000 440.590 1500.000 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 321.680 1500.000 322.280 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 1496.000 534.430 1500.000 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 1496.000 553.290 1500.000 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 1496.000 609.410 1500.000 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 1496.000 628.270 1500.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 461.080 1500.000 461.680 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 496.440 1500.000 497.040 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 513.440 1500.000 514.040 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 1496.000 684.390 1500.000 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 565.800 1500.000 566.400 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 112.240 1500.000 112.840 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 1496.000 252.910 1500.000 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 1496.000 290.630 1500.000 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 1496.000 84.550 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 1496.000 121.810 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 8.200 1500.000 8.800 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 1496.000 102.950 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 234.640 1500.000 235.240 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 304.680 1500.000 305.280 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 339.360 1500.000 339.960 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 25.200 1500.000 25.800 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 1496.000 234.510 1500.000 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 129.920 1500.000 130.520 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 164.600 1500.000 165.200 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1225.400 4.000 1226.000 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1260.760 4.000 1261.360 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1246.480 1500.000 1247.080 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.810 1496.000 1303.090 1500.000 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.670 1496.000 1321.950 1500.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1298.840 1500.000 1299.440 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1278.440 4.000 1279.040 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 1496.000 1359.210 1500.000 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.790 1496.000 1378.070 1500.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.890 0.000 1371.170 4.000 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 182.280 1500.000 182.880 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1333.520 1500.000 1334.120 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1351.200 1500.000 1351.800 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1313.800 4.000 1314.400 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.510 1496.000 1415.790 1500.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.250 0.000 1401.530 4.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 1496.000 1471.910 1500.000 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1331.480 4.000 1332.080 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.160 4.000 1349.760 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1420.560 1500.000 1421.160 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.840 4.000 1367.440 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.790 0.000 1447.070 4.000 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1402.200 4.000 1402.800 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 0.000 1462.250 4.000 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.150 0.000 1477.430 4.000 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1455.920 1500.000 1456.520 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1437.560 4.000 1438.160 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1490.600 1500.000 1491.200 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1490.600 4.000 1491.200 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 1496.000 365.610 1500.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 269.320 1500.000 269.920 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 287.000 1500.000 287.600 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 1496.000 496.710 1500.000 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 42.880 1500.000 43.480 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 374.040 1500.000 374.640 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 1496.000 571.690 1500.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 426.400 1500.000 427.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 478.760 1500.000 479.360 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 548.800 1500.000 549.400 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 583.480 1500.000 584.080 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 766.400 4.000 767.000 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.760 4.000 802.360 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1496.000 721.650 1500.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 635.840 1500.000 636.440 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 1496.000 740.510 1500.000 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.120 4.000 837.720 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 1496.000 177.930 1500.000 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 653.520 1500.000 654.120 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.800 4.000 855.400 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 0.000 825.610 4.000 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 722.880 1500.000 723.480 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 1496.000 797.090 1500.000 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 872.480 4.000 873.080 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 1496.000 196.790 1500.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.160 4.000 890.760 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 0.000 931.870 4.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 740.560 1500.000 741.160 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 1496.000 890.470 1500.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 0.000 977.410 4.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 0.000 992.590 4.000 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 775.240 1500.000 775.840 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 0.000 1022.490 4.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 95.240 1500.000 95.840 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 1496.000 928.190 1500.000 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 809.920 1500.000 810.520 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 827.600 1500.000 828.200 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.200 4.000 943.800 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 978.560 4.000 979.160 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 1496.000 965.450 1500.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 1496.000 984.310 1500.000 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 0.000 1128.750 4.000 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 862.280 1500.000 862.880 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.750 1496.000 1022.030 1500.000 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.280 4.000 1049.880 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.960 4.000 1067.560 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 879.960 1500.000 880.560 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 897.640 1500.000 898.240 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.870 1496.000 1078.150 1500.000 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 0.000 1174.290 4.000 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 932.320 1500.000 932.920 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.000 4.000 1120.600 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 950.000 1500.000 950.600 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.730 1496.000 1097.010 1500.000 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 967.000 1500.000 967.600 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 0.000 1219.830 4.000 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1234.730 0.000 1235.010 4.000 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 0.000 1250.190 4.000 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1019.360 1500.000 1019.960 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1054.720 1500.000 1055.320 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1071.720 1500.000 1072.320 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1107.080 1500.000 1107.680 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.570 1496.000 1190.850 1500.000 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1141.760 1500.000 1142.360 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.810 0.000 1280.090 4.000 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1158.760 1500.000 1159.360 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.990 0.000 1295.270 4.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.830 1496.000 1228.110 1500.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1211.120 1500.000 1211.720 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 1496.000 1265.830 1500.000 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.720 4.000 1208.320 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 1496.000 309.490 1500.000 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 1496.000 46.830 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 1496.000 65.690 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 252.320 1500.000 252.920 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 1496.000 384.470 1500.000 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 1496.000 459.450 1500.000 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 1496.000 478.310 1500.000 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 357.040 1500.000 357.640 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 408.720 1500.000 409.320 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 1496.000 646.670 1500.000 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 531.120 1500.000 531.720 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 59.880 1500.000 60.480 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 147.600 1500.000 148.200 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 1496.000 327.890 1500.000 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 1496.000 27.970 1500.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 7.225 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.080 1489.500 ;
      LAYER met2 ;
        RECT 6.990 1495.720 9.010 1496.410 ;
        RECT 9.850 1495.720 27.410 1496.410 ;
        RECT 28.250 1495.720 46.270 1496.410 ;
        RECT 47.110 1495.720 65.130 1496.410 ;
        RECT 65.970 1495.720 83.990 1496.410 ;
        RECT 84.830 1495.720 102.390 1496.410 ;
        RECT 103.230 1495.720 121.250 1496.410 ;
        RECT 122.090 1495.720 140.110 1496.410 ;
        RECT 140.950 1495.720 158.970 1496.410 ;
        RECT 159.810 1495.720 177.370 1496.410 ;
        RECT 178.210 1495.720 196.230 1496.410 ;
        RECT 197.070 1495.720 215.090 1496.410 ;
        RECT 215.930 1495.720 233.950 1496.410 ;
        RECT 234.790 1495.720 252.350 1496.410 ;
        RECT 253.190 1495.720 271.210 1496.410 ;
        RECT 272.050 1495.720 290.070 1496.410 ;
        RECT 290.910 1495.720 308.930 1496.410 ;
        RECT 309.770 1495.720 327.330 1496.410 ;
        RECT 328.170 1495.720 346.190 1496.410 ;
        RECT 347.030 1495.720 365.050 1496.410 ;
        RECT 365.890 1495.720 383.910 1496.410 ;
        RECT 384.750 1495.720 402.770 1496.410 ;
        RECT 403.610 1495.720 421.170 1496.410 ;
        RECT 422.010 1495.720 440.030 1496.410 ;
        RECT 440.870 1495.720 458.890 1496.410 ;
        RECT 459.730 1495.720 477.750 1496.410 ;
        RECT 478.590 1495.720 496.150 1496.410 ;
        RECT 496.990 1495.720 515.010 1496.410 ;
        RECT 515.850 1495.720 533.870 1496.410 ;
        RECT 534.710 1495.720 552.730 1496.410 ;
        RECT 553.570 1495.720 571.130 1496.410 ;
        RECT 571.970 1495.720 589.990 1496.410 ;
        RECT 590.830 1495.720 608.850 1496.410 ;
        RECT 609.690 1495.720 627.710 1496.410 ;
        RECT 628.550 1495.720 646.110 1496.410 ;
        RECT 646.950 1495.720 664.970 1496.410 ;
        RECT 665.810 1495.720 683.830 1496.410 ;
        RECT 684.670 1495.720 702.690 1496.410 ;
        RECT 703.530 1495.720 721.090 1496.410 ;
        RECT 721.930 1495.720 739.950 1496.410 ;
        RECT 740.790 1495.720 758.810 1496.410 ;
        RECT 759.650 1495.720 777.670 1496.410 ;
        RECT 778.510 1495.720 796.530 1496.410 ;
        RECT 797.370 1495.720 814.930 1496.410 ;
        RECT 815.770 1495.720 833.790 1496.410 ;
        RECT 834.630 1495.720 852.650 1496.410 ;
        RECT 853.490 1495.720 871.510 1496.410 ;
        RECT 872.350 1495.720 889.910 1496.410 ;
        RECT 890.750 1495.720 908.770 1496.410 ;
        RECT 909.610 1495.720 927.630 1496.410 ;
        RECT 928.470 1495.720 946.490 1496.410 ;
        RECT 947.330 1495.720 964.890 1496.410 ;
        RECT 965.730 1495.720 983.750 1496.410 ;
        RECT 984.590 1495.720 1002.610 1496.410 ;
        RECT 1003.450 1495.720 1021.470 1496.410 ;
        RECT 1022.310 1495.720 1039.870 1496.410 ;
        RECT 1040.710 1495.720 1058.730 1496.410 ;
        RECT 1059.570 1495.720 1077.590 1496.410 ;
        RECT 1078.430 1495.720 1096.450 1496.410 ;
        RECT 1097.290 1495.720 1114.850 1496.410 ;
        RECT 1115.690 1495.720 1133.710 1496.410 ;
        RECT 1134.550 1495.720 1152.570 1496.410 ;
        RECT 1153.410 1495.720 1171.430 1496.410 ;
        RECT 1172.270 1495.720 1190.290 1496.410 ;
        RECT 1191.130 1495.720 1208.690 1496.410 ;
        RECT 1209.530 1495.720 1227.550 1496.410 ;
        RECT 1228.390 1495.720 1246.410 1496.410 ;
        RECT 1247.250 1495.720 1265.270 1496.410 ;
        RECT 1266.110 1495.720 1283.670 1496.410 ;
        RECT 1284.510 1495.720 1302.530 1496.410 ;
        RECT 1303.370 1495.720 1321.390 1496.410 ;
        RECT 1322.230 1495.720 1340.250 1496.410 ;
        RECT 1341.090 1495.720 1358.650 1496.410 ;
        RECT 1359.490 1495.720 1377.510 1496.410 ;
        RECT 1378.350 1495.720 1396.370 1496.410 ;
        RECT 1397.210 1495.720 1415.230 1496.410 ;
        RECT 1416.070 1495.720 1433.630 1496.410 ;
        RECT 1434.470 1495.720 1452.490 1496.410 ;
        RECT 1453.330 1495.720 1471.350 1496.410 ;
        RECT 1472.190 1495.720 1490.210 1496.410 ;
        RECT 1491.050 1495.720 1492.600 1496.410 ;
        RECT 6.990 4.280 1492.600 1495.720 ;
        RECT 6.990 3.670 7.170 4.280 ;
        RECT 8.010 3.670 21.890 4.280 ;
        RECT 22.730 3.670 37.070 4.280 ;
        RECT 37.910 3.670 52.250 4.280 ;
        RECT 53.090 3.670 67.430 4.280 ;
        RECT 68.270 3.670 82.610 4.280 ;
        RECT 83.450 3.670 97.790 4.280 ;
        RECT 98.630 3.670 112.970 4.280 ;
        RECT 113.810 3.670 128.150 4.280 ;
        RECT 128.990 3.670 143.330 4.280 ;
        RECT 144.170 3.670 158.510 4.280 ;
        RECT 159.350 3.670 173.690 4.280 ;
        RECT 174.530 3.670 188.870 4.280 ;
        RECT 189.710 3.670 204.050 4.280 ;
        RECT 204.890 3.670 219.230 4.280 ;
        RECT 220.070 3.670 234.410 4.280 ;
        RECT 235.250 3.670 249.590 4.280 ;
        RECT 250.430 3.670 264.310 4.280 ;
        RECT 265.150 3.670 279.490 4.280 ;
        RECT 280.330 3.670 294.670 4.280 ;
        RECT 295.510 3.670 309.850 4.280 ;
        RECT 310.690 3.670 325.030 4.280 ;
        RECT 325.870 3.670 340.210 4.280 ;
        RECT 341.050 3.670 355.390 4.280 ;
        RECT 356.230 3.670 370.570 4.280 ;
        RECT 371.410 3.670 385.750 4.280 ;
        RECT 386.590 3.670 400.930 4.280 ;
        RECT 401.770 3.670 416.110 4.280 ;
        RECT 416.950 3.670 431.290 4.280 ;
        RECT 432.130 3.670 446.470 4.280 ;
        RECT 447.310 3.670 461.650 4.280 ;
        RECT 462.490 3.670 476.830 4.280 ;
        RECT 477.670 3.670 492.010 4.280 ;
        RECT 492.850 3.670 507.190 4.280 ;
        RECT 508.030 3.670 521.910 4.280 ;
        RECT 522.750 3.670 537.090 4.280 ;
        RECT 537.930 3.670 552.270 4.280 ;
        RECT 553.110 3.670 567.450 4.280 ;
        RECT 568.290 3.670 582.630 4.280 ;
        RECT 583.470 3.670 597.810 4.280 ;
        RECT 598.650 3.670 612.990 4.280 ;
        RECT 613.830 3.670 628.170 4.280 ;
        RECT 629.010 3.670 643.350 4.280 ;
        RECT 644.190 3.670 658.530 4.280 ;
        RECT 659.370 3.670 673.710 4.280 ;
        RECT 674.550 3.670 688.890 4.280 ;
        RECT 689.730 3.670 704.070 4.280 ;
        RECT 704.910 3.670 719.250 4.280 ;
        RECT 720.090 3.670 734.430 4.280 ;
        RECT 735.270 3.670 749.610 4.280 ;
        RECT 750.450 3.670 764.330 4.280 ;
        RECT 765.170 3.670 779.510 4.280 ;
        RECT 780.350 3.670 794.690 4.280 ;
        RECT 795.530 3.670 809.870 4.280 ;
        RECT 810.710 3.670 825.050 4.280 ;
        RECT 825.890 3.670 840.230 4.280 ;
        RECT 841.070 3.670 855.410 4.280 ;
        RECT 856.250 3.670 870.590 4.280 ;
        RECT 871.430 3.670 885.770 4.280 ;
        RECT 886.610 3.670 900.950 4.280 ;
        RECT 901.790 3.670 916.130 4.280 ;
        RECT 916.970 3.670 931.310 4.280 ;
        RECT 932.150 3.670 946.490 4.280 ;
        RECT 947.330 3.670 961.670 4.280 ;
        RECT 962.510 3.670 976.850 4.280 ;
        RECT 977.690 3.670 992.030 4.280 ;
        RECT 992.870 3.670 1007.210 4.280 ;
        RECT 1008.050 3.670 1021.930 4.280 ;
        RECT 1022.770 3.670 1037.110 4.280 ;
        RECT 1037.950 3.670 1052.290 4.280 ;
        RECT 1053.130 3.670 1067.470 4.280 ;
        RECT 1068.310 3.670 1082.650 4.280 ;
        RECT 1083.490 3.670 1097.830 4.280 ;
        RECT 1098.670 3.670 1113.010 4.280 ;
        RECT 1113.850 3.670 1128.190 4.280 ;
        RECT 1129.030 3.670 1143.370 4.280 ;
        RECT 1144.210 3.670 1158.550 4.280 ;
        RECT 1159.390 3.670 1173.730 4.280 ;
        RECT 1174.570 3.670 1188.910 4.280 ;
        RECT 1189.750 3.670 1204.090 4.280 ;
        RECT 1204.930 3.670 1219.270 4.280 ;
        RECT 1220.110 3.670 1234.450 4.280 ;
        RECT 1235.290 3.670 1249.630 4.280 ;
        RECT 1250.470 3.670 1264.350 4.280 ;
        RECT 1265.190 3.670 1279.530 4.280 ;
        RECT 1280.370 3.670 1294.710 4.280 ;
        RECT 1295.550 3.670 1309.890 4.280 ;
        RECT 1310.730 3.670 1325.070 4.280 ;
        RECT 1325.910 3.670 1340.250 4.280 ;
        RECT 1341.090 3.670 1355.430 4.280 ;
        RECT 1356.270 3.670 1370.610 4.280 ;
        RECT 1371.450 3.670 1385.790 4.280 ;
        RECT 1386.630 3.670 1400.970 4.280 ;
        RECT 1401.810 3.670 1416.150 4.280 ;
        RECT 1416.990 3.670 1431.330 4.280 ;
        RECT 1432.170 3.670 1446.510 4.280 ;
        RECT 1447.350 3.670 1461.690 4.280 ;
        RECT 1462.530 3.670 1476.870 4.280 ;
        RECT 1477.710 3.670 1492.050 4.280 ;
      LAYER met3 ;
        RECT 4.400 1490.200 1495.600 1491.065 ;
        RECT 4.000 1473.920 1496.000 1490.200 ;
        RECT 4.400 1472.520 1495.600 1473.920 ;
        RECT 4.000 1456.920 1496.000 1472.520 ;
        RECT 4.000 1456.240 1495.600 1456.920 ;
        RECT 4.400 1455.520 1495.600 1456.240 ;
        RECT 4.400 1454.840 1496.000 1455.520 ;
        RECT 4.000 1439.240 1496.000 1454.840 ;
        RECT 4.000 1438.560 1495.600 1439.240 ;
        RECT 4.400 1437.840 1495.600 1438.560 ;
        RECT 4.400 1437.160 1496.000 1437.840 ;
        RECT 4.000 1421.560 1496.000 1437.160 ;
        RECT 4.000 1420.880 1495.600 1421.560 ;
        RECT 4.400 1420.160 1495.600 1420.880 ;
        RECT 4.400 1419.480 1496.000 1420.160 ;
        RECT 4.000 1404.560 1496.000 1419.480 ;
        RECT 4.000 1403.200 1495.600 1404.560 ;
        RECT 4.400 1403.160 1495.600 1403.200 ;
        RECT 4.400 1401.800 1496.000 1403.160 ;
        RECT 4.000 1386.880 1496.000 1401.800 ;
        RECT 4.000 1385.520 1495.600 1386.880 ;
        RECT 4.400 1385.480 1495.600 1385.520 ;
        RECT 4.400 1384.120 1496.000 1385.480 ;
        RECT 4.000 1369.200 1496.000 1384.120 ;
        RECT 4.000 1367.840 1495.600 1369.200 ;
        RECT 4.400 1367.800 1495.600 1367.840 ;
        RECT 4.400 1366.440 1496.000 1367.800 ;
        RECT 4.000 1352.200 1496.000 1366.440 ;
        RECT 4.000 1350.800 1495.600 1352.200 ;
        RECT 4.000 1350.160 1496.000 1350.800 ;
        RECT 4.400 1348.760 1496.000 1350.160 ;
        RECT 4.000 1334.520 1496.000 1348.760 ;
        RECT 4.000 1333.120 1495.600 1334.520 ;
        RECT 4.000 1332.480 1496.000 1333.120 ;
        RECT 4.400 1331.080 1496.000 1332.480 ;
        RECT 4.000 1316.840 1496.000 1331.080 ;
        RECT 4.000 1315.440 1495.600 1316.840 ;
        RECT 4.000 1314.800 1496.000 1315.440 ;
        RECT 4.400 1313.400 1496.000 1314.800 ;
        RECT 4.000 1299.840 1496.000 1313.400 ;
        RECT 4.000 1298.440 1495.600 1299.840 ;
        RECT 4.000 1297.120 1496.000 1298.440 ;
        RECT 4.400 1295.720 1496.000 1297.120 ;
        RECT 4.000 1282.160 1496.000 1295.720 ;
        RECT 4.000 1280.760 1495.600 1282.160 ;
        RECT 4.000 1279.440 1496.000 1280.760 ;
        RECT 4.400 1278.040 1496.000 1279.440 ;
        RECT 4.000 1264.480 1496.000 1278.040 ;
        RECT 4.000 1263.080 1495.600 1264.480 ;
        RECT 4.000 1261.760 1496.000 1263.080 ;
        RECT 4.400 1260.360 1496.000 1261.760 ;
        RECT 4.000 1247.480 1496.000 1260.360 ;
        RECT 4.000 1246.080 1495.600 1247.480 ;
        RECT 4.000 1244.080 1496.000 1246.080 ;
        RECT 4.400 1242.680 1496.000 1244.080 ;
        RECT 4.000 1229.800 1496.000 1242.680 ;
        RECT 4.000 1228.400 1495.600 1229.800 ;
        RECT 4.000 1226.400 1496.000 1228.400 ;
        RECT 4.400 1225.000 1496.000 1226.400 ;
        RECT 4.000 1212.120 1496.000 1225.000 ;
        RECT 4.000 1210.720 1495.600 1212.120 ;
        RECT 4.000 1208.720 1496.000 1210.720 ;
        RECT 4.400 1207.320 1496.000 1208.720 ;
        RECT 4.000 1195.120 1496.000 1207.320 ;
        RECT 4.000 1193.720 1495.600 1195.120 ;
        RECT 4.000 1191.040 1496.000 1193.720 ;
        RECT 4.400 1189.640 1496.000 1191.040 ;
        RECT 4.000 1177.440 1496.000 1189.640 ;
        RECT 4.000 1176.040 1495.600 1177.440 ;
        RECT 4.000 1173.360 1496.000 1176.040 ;
        RECT 4.400 1171.960 1496.000 1173.360 ;
        RECT 4.000 1159.760 1496.000 1171.960 ;
        RECT 4.000 1158.360 1495.600 1159.760 ;
        RECT 4.000 1155.680 1496.000 1158.360 ;
        RECT 4.400 1154.280 1496.000 1155.680 ;
        RECT 4.000 1142.760 1496.000 1154.280 ;
        RECT 4.000 1141.360 1495.600 1142.760 ;
        RECT 4.000 1138.000 1496.000 1141.360 ;
        RECT 4.400 1136.600 1496.000 1138.000 ;
        RECT 4.000 1125.080 1496.000 1136.600 ;
        RECT 4.000 1123.680 1495.600 1125.080 ;
        RECT 4.000 1121.000 1496.000 1123.680 ;
        RECT 4.400 1119.600 1496.000 1121.000 ;
        RECT 4.000 1108.080 1496.000 1119.600 ;
        RECT 4.000 1106.680 1495.600 1108.080 ;
        RECT 4.000 1103.320 1496.000 1106.680 ;
        RECT 4.400 1101.920 1496.000 1103.320 ;
        RECT 4.000 1090.400 1496.000 1101.920 ;
        RECT 4.000 1089.000 1495.600 1090.400 ;
        RECT 4.000 1085.640 1496.000 1089.000 ;
        RECT 4.400 1084.240 1496.000 1085.640 ;
        RECT 4.000 1072.720 1496.000 1084.240 ;
        RECT 4.000 1071.320 1495.600 1072.720 ;
        RECT 4.000 1067.960 1496.000 1071.320 ;
        RECT 4.400 1066.560 1496.000 1067.960 ;
        RECT 4.000 1055.720 1496.000 1066.560 ;
        RECT 4.000 1054.320 1495.600 1055.720 ;
        RECT 4.000 1050.280 1496.000 1054.320 ;
        RECT 4.400 1048.880 1496.000 1050.280 ;
        RECT 4.000 1038.040 1496.000 1048.880 ;
        RECT 4.000 1036.640 1495.600 1038.040 ;
        RECT 4.000 1032.600 1496.000 1036.640 ;
        RECT 4.400 1031.200 1496.000 1032.600 ;
        RECT 4.000 1020.360 1496.000 1031.200 ;
        RECT 4.000 1018.960 1495.600 1020.360 ;
        RECT 4.000 1014.920 1496.000 1018.960 ;
        RECT 4.400 1013.520 1496.000 1014.920 ;
        RECT 4.000 1003.360 1496.000 1013.520 ;
        RECT 4.000 1001.960 1495.600 1003.360 ;
        RECT 4.000 997.240 1496.000 1001.960 ;
        RECT 4.400 995.840 1496.000 997.240 ;
        RECT 4.000 985.680 1496.000 995.840 ;
        RECT 4.000 984.280 1495.600 985.680 ;
        RECT 4.000 979.560 1496.000 984.280 ;
        RECT 4.400 978.160 1496.000 979.560 ;
        RECT 4.000 968.000 1496.000 978.160 ;
        RECT 4.000 966.600 1495.600 968.000 ;
        RECT 4.000 961.880 1496.000 966.600 ;
        RECT 4.400 960.480 1496.000 961.880 ;
        RECT 4.000 951.000 1496.000 960.480 ;
        RECT 4.000 949.600 1495.600 951.000 ;
        RECT 4.000 944.200 1496.000 949.600 ;
        RECT 4.400 942.800 1496.000 944.200 ;
        RECT 4.000 933.320 1496.000 942.800 ;
        RECT 4.000 931.920 1495.600 933.320 ;
        RECT 4.000 926.520 1496.000 931.920 ;
        RECT 4.400 925.120 1496.000 926.520 ;
        RECT 4.000 915.640 1496.000 925.120 ;
        RECT 4.000 914.240 1495.600 915.640 ;
        RECT 4.000 908.840 1496.000 914.240 ;
        RECT 4.400 907.440 1496.000 908.840 ;
        RECT 4.000 898.640 1496.000 907.440 ;
        RECT 4.000 897.240 1495.600 898.640 ;
        RECT 4.000 891.160 1496.000 897.240 ;
        RECT 4.400 889.760 1496.000 891.160 ;
        RECT 4.000 880.960 1496.000 889.760 ;
        RECT 4.000 879.560 1495.600 880.960 ;
        RECT 4.000 873.480 1496.000 879.560 ;
        RECT 4.400 872.080 1496.000 873.480 ;
        RECT 4.000 863.280 1496.000 872.080 ;
        RECT 4.000 861.880 1495.600 863.280 ;
        RECT 4.000 855.800 1496.000 861.880 ;
        RECT 4.400 854.400 1496.000 855.800 ;
        RECT 4.000 846.280 1496.000 854.400 ;
        RECT 4.000 844.880 1495.600 846.280 ;
        RECT 4.000 838.120 1496.000 844.880 ;
        RECT 4.400 836.720 1496.000 838.120 ;
        RECT 4.000 828.600 1496.000 836.720 ;
        RECT 4.000 827.200 1495.600 828.600 ;
        RECT 4.000 820.440 1496.000 827.200 ;
        RECT 4.400 819.040 1496.000 820.440 ;
        RECT 4.000 810.920 1496.000 819.040 ;
        RECT 4.000 809.520 1495.600 810.920 ;
        RECT 4.000 802.760 1496.000 809.520 ;
        RECT 4.400 801.360 1496.000 802.760 ;
        RECT 4.000 793.920 1496.000 801.360 ;
        RECT 4.000 792.520 1495.600 793.920 ;
        RECT 4.000 785.080 1496.000 792.520 ;
        RECT 4.400 783.680 1496.000 785.080 ;
        RECT 4.000 776.240 1496.000 783.680 ;
        RECT 4.000 774.840 1495.600 776.240 ;
        RECT 4.000 767.400 1496.000 774.840 ;
        RECT 4.400 766.000 1496.000 767.400 ;
        RECT 4.000 759.240 1496.000 766.000 ;
        RECT 4.000 757.840 1495.600 759.240 ;
        RECT 4.000 750.400 1496.000 757.840 ;
        RECT 4.400 749.000 1496.000 750.400 ;
        RECT 4.000 741.560 1496.000 749.000 ;
        RECT 4.000 740.160 1495.600 741.560 ;
        RECT 4.000 732.720 1496.000 740.160 ;
        RECT 4.400 731.320 1496.000 732.720 ;
        RECT 4.000 723.880 1496.000 731.320 ;
        RECT 4.000 722.480 1495.600 723.880 ;
        RECT 4.000 715.040 1496.000 722.480 ;
        RECT 4.400 713.640 1496.000 715.040 ;
        RECT 4.000 706.880 1496.000 713.640 ;
        RECT 4.000 705.480 1495.600 706.880 ;
        RECT 4.000 697.360 1496.000 705.480 ;
        RECT 4.400 695.960 1496.000 697.360 ;
        RECT 4.000 689.200 1496.000 695.960 ;
        RECT 4.000 687.800 1495.600 689.200 ;
        RECT 4.000 679.680 1496.000 687.800 ;
        RECT 4.400 678.280 1496.000 679.680 ;
        RECT 4.000 671.520 1496.000 678.280 ;
        RECT 4.000 670.120 1495.600 671.520 ;
        RECT 4.000 662.000 1496.000 670.120 ;
        RECT 4.400 660.600 1496.000 662.000 ;
        RECT 4.000 654.520 1496.000 660.600 ;
        RECT 4.000 653.120 1495.600 654.520 ;
        RECT 4.000 644.320 1496.000 653.120 ;
        RECT 4.400 642.920 1496.000 644.320 ;
        RECT 4.000 636.840 1496.000 642.920 ;
        RECT 4.000 635.440 1495.600 636.840 ;
        RECT 4.000 626.640 1496.000 635.440 ;
        RECT 4.400 625.240 1496.000 626.640 ;
        RECT 4.000 619.160 1496.000 625.240 ;
        RECT 4.000 617.760 1495.600 619.160 ;
        RECT 4.000 608.960 1496.000 617.760 ;
        RECT 4.400 607.560 1496.000 608.960 ;
        RECT 4.000 602.160 1496.000 607.560 ;
        RECT 4.000 600.760 1495.600 602.160 ;
        RECT 4.000 591.280 1496.000 600.760 ;
        RECT 4.400 589.880 1496.000 591.280 ;
        RECT 4.000 584.480 1496.000 589.880 ;
        RECT 4.000 583.080 1495.600 584.480 ;
        RECT 4.000 573.600 1496.000 583.080 ;
        RECT 4.400 572.200 1496.000 573.600 ;
        RECT 4.000 566.800 1496.000 572.200 ;
        RECT 4.000 565.400 1495.600 566.800 ;
        RECT 4.000 555.920 1496.000 565.400 ;
        RECT 4.400 554.520 1496.000 555.920 ;
        RECT 4.000 549.800 1496.000 554.520 ;
        RECT 4.000 548.400 1495.600 549.800 ;
        RECT 4.000 538.240 1496.000 548.400 ;
        RECT 4.400 536.840 1496.000 538.240 ;
        RECT 4.000 532.120 1496.000 536.840 ;
        RECT 4.000 530.720 1495.600 532.120 ;
        RECT 4.000 520.560 1496.000 530.720 ;
        RECT 4.400 519.160 1496.000 520.560 ;
        RECT 4.000 514.440 1496.000 519.160 ;
        RECT 4.000 513.040 1495.600 514.440 ;
        RECT 4.000 502.880 1496.000 513.040 ;
        RECT 4.400 501.480 1496.000 502.880 ;
        RECT 4.000 497.440 1496.000 501.480 ;
        RECT 4.000 496.040 1495.600 497.440 ;
        RECT 4.000 485.200 1496.000 496.040 ;
        RECT 4.400 483.800 1496.000 485.200 ;
        RECT 4.000 479.760 1496.000 483.800 ;
        RECT 4.000 478.360 1495.600 479.760 ;
        RECT 4.000 467.520 1496.000 478.360 ;
        RECT 4.400 466.120 1496.000 467.520 ;
        RECT 4.000 462.080 1496.000 466.120 ;
        RECT 4.000 460.680 1495.600 462.080 ;
        RECT 4.000 449.840 1496.000 460.680 ;
        RECT 4.400 448.440 1496.000 449.840 ;
        RECT 4.000 445.080 1496.000 448.440 ;
        RECT 4.000 443.680 1495.600 445.080 ;
        RECT 4.000 432.160 1496.000 443.680 ;
        RECT 4.400 430.760 1496.000 432.160 ;
        RECT 4.000 427.400 1496.000 430.760 ;
        RECT 4.000 426.000 1495.600 427.400 ;
        RECT 4.000 414.480 1496.000 426.000 ;
        RECT 4.400 413.080 1496.000 414.480 ;
        RECT 4.000 409.720 1496.000 413.080 ;
        RECT 4.000 408.320 1495.600 409.720 ;
        RECT 4.000 396.800 1496.000 408.320 ;
        RECT 4.400 395.400 1496.000 396.800 ;
        RECT 4.000 392.720 1496.000 395.400 ;
        RECT 4.000 391.320 1495.600 392.720 ;
        RECT 4.000 379.800 1496.000 391.320 ;
        RECT 4.400 378.400 1496.000 379.800 ;
        RECT 4.000 375.040 1496.000 378.400 ;
        RECT 4.000 373.640 1495.600 375.040 ;
        RECT 4.000 362.120 1496.000 373.640 ;
        RECT 4.400 360.720 1496.000 362.120 ;
        RECT 4.000 358.040 1496.000 360.720 ;
        RECT 4.000 356.640 1495.600 358.040 ;
        RECT 4.000 344.440 1496.000 356.640 ;
        RECT 4.400 343.040 1496.000 344.440 ;
        RECT 4.000 340.360 1496.000 343.040 ;
        RECT 4.000 338.960 1495.600 340.360 ;
        RECT 4.000 326.760 1496.000 338.960 ;
        RECT 4.400 325.360 1496.000 326.760 ;
        RECT 4.000 322.680 1496.000 325.360 ;
        RECT 4.000 321.280 1495.600 322.680 ;
        RECT 4.000 309.080 1496.000 321.280 ;
        RECT 4.400 307.680 1496.000 309.080 ;
        RECT 4.000 305.680 1496.000 307.680 ;
        RECT 4.000 304.280 1495.600 305.680 ;
        RECT 4.000 291.400 1496.000 304.280 ;
        RECT 4.400 290.000 1496.000 291.400 ;
        RECT 4.000 288.000 1496.000 290.000 ;
        RECT 4.000 286.600 1495.600 288.000 ;
        RECT 4.000 273.720 1496.000 286.600 ;
        RECT 4.400 272.320 1496.000 273.720 ;
        RECT 4.000 270.320 1496.000 272.320 ;
        RECT 4.000 268.920 1495.600 270.320 ;
        RECT 4.000 256.040 1496.000 268.920 ;
        RECT 4.400 254.640 1496.000 256.040 ;
        RECT 4.000 253.320 1496.000 254.640 ;
        RECT 4.000 251.920 1495.600 253.320 ;
        RECT 4.000 238.360 1496.000 251.920 ;
        RECT 4.400 236.960 1496.000 238.360 ;
        RECT 4.000 235.640 1496.000 236.960 ;
        RECT 4.000 234.240 1495.600 235.640 ;
        RECT 4.000 220.680 1496.000 234.240 ;
        RECT 4.400 219.280 1496.000 220.680 ;
        RECT 4.000 217.960 1496.000 219.280 ;
        RECT 4.000 216.560 1495.600 217.960 ;
        RECT 4.000 203.000 1496.000 216.560 ;
        RECT 4.400 201.600 1496.000 203.000 ;
        RECT 4.000 200.960 1496.000 201.600 ;
        RECT 4.000 199.560 1495.600 200.960 ;
        RECT 4.000 185.320 1496.000 199.560 ;
        RECT 4.400 183.920 1496.000 185.320 ;
        RECT 4.000 183.280 1496.000 183.920 ;
        RECT 4.000 181.880 1495.600 183.280 ;
        RECT 4.000 167.640 1496.000 181.880 ;
        RECT 4.400 166.240 1496.000 167.640 ;
        RECT 4.000 165.600 1496.000 166.240 ;
        RECT 4.000 164.200 1495.600 165.600 ;
        RECT 4.000 149.960 1496.000 164.200 ;
        RECT 4.400 148.600 1496.000 149.960 ;
        RECT 4.400 148.560 1495.600 148.600 ;
        RECT 4.000 147.200 1495.600 148.560 ;
        RECT 4.000 132.280 1496.000 147.200 ;
        RECT 4.400 130.920 1496.000 132.280 ;
        RECT 4.400 130.880 1495.600 130.920 ;
        RECT 4.000 129.520 1495.600 130.880 ;
        RECT 4.000 114.600 1496.000 129.520 ;
        RECT 4.400 113.240 1496.000 114.600 ;
        RECT 4.400 113.200 1495.600 113.240 ;
        RECT 4.000 111.840 1495.600 113.200 ;
        RECT 4.000 96.920 1496.000 111.840 ;
        RECT 4.400 96.240 1496.000 96.920 ;
        RECT 4.400 95.520 1495.600 96.240 ;
        RECT 4.000 94.840 1495.600 95.520 ;
        RECT 4.000 79.240 1496.000 94.840 ;
        RECT 4.400 78.560 1496.000 79.240 ;
        RECT 4.400 77.840 1495.600 78.560 ;
        RECT 4.000 77.160 1495.600 77.840 ;
        RECT 4.000 61.560 1496.000 77.160 ;
        RECT 4.400 60.880 1496.000 61.560 ;
        RECT 4.400 60.160 1495.600 60.880 ;
        RECT 4.000 59.480 1495.600 60.160 ;
        RECT 4.000 43.880 1496.000 59.480 ;
        RECT 4.400 42.480 1495.600 43.880 ;
        RECT 4.000 26.200 1496.000 42.480 ;
        RECT 4.400 24.800 1495.600 26.200 ;
        RECT 4.000 9.200 1496.000 24.800 ;
        RECT 4.400 8.335 1495.600 9.200 ;
      LAYER met4 ;
        RECT 100.575 11.735 174.240 1486.305 ;
        RECT 176.640 11.735 251.040 1486.305 ;
        RECT 253.440 11.735 327.840 1486.305 ;
        RECT 330.240 11.735 404.640 1486.305 ;
        RECT 407.040 11.735 481.440 1486.305 ;
        RECT 483.840 11.735 558.240 1486.305 ;
        RECT 560.640 11.735 635.040 1486.305 ;
        RECT 637.440 11.735 711.840 1486.305 ;
        RECT 714.240 11.735 788.640 1486.305 ;
        RECT 791.040 11.735 865.440 1486.305 ;
        RECT 867.840 11.735 942.240 1486.305 ;
        RECT 944.640 11.735 1019.040 1486.305 ;
        RECT 1021.440 11.735 1095.840 1486.305 ;
        RECT 1098.240 11.735 1110.145 1486.305 ;
  END
END core
END LIBRARY

