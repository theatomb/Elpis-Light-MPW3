VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO io_output_arbiter
  CLASS BLOCK ;
  FOREIGN io_output_arbiter ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 75.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END clk
  PIN data_core0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END data_core0[0]
  PIN data_core0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END data_core0[10]
  PIN data_core0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END data_core0[11]
  PIN data_core0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END data_core0[12]
  PIN data_core0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 71.000 22.910 75.000 ;
    END
  END data_core0[13]
  PIN data_core0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END data_core0[14]
  PIN data_core0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 71.000 31.190 75.000 ;
    END
  END data_core0[15]
  PIN data_core0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 34.040 75.000 34.640 ;
    END
  END data_core0[16]
  PIN data_core0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END data_core0[17]
  PIN data_core0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 44.240 75.000 44.840 ;
    END
  END data_core0[18]
  PIN data_core0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 71.000 35.330 75.000 ;
    END
  END data_core0[19]
  PIN data_core0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 2.080 75.000 2.680 ;
    END
  END data_core0[1]
  PIN data_core0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END data_core0[20]
  PIN data_core0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 49.680 75.000 50.280 ;
    END
  END data_core0[21]
  PIN data_core0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 71.000 47.750 75.000 ;
    END
  END data_core0[22]
  PIN data_core0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END data_core0[23]
  PIN data_core0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END data_core0[24]
  PIN data_core0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END data_core0[25]
  PIN data_core0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 60.560 75.000 61.160 ;
    END
  END data_core0[26]
  PIN data_core0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END data_core0[27]
  PIN data_core0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END data_core0[28]
  PIN data_core0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 71.000 64.310 75.000 ;
    END
  END data_core0[29]
  PIN data_core0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 71.000 2.210 75.000 ;
    END
  END data_core0[2]
  PIN data_core0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 71.440 75.000 72.040 ;
    END
  END data_core0[30]
  PIN data_core0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 71.000 72.590 75.000 ;
    END
  END data_core0[31]
  PIN data_core0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 71.000 6.350 75.000 ;
    END
  END data_core0[3]
  PIN data_core0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END data_core0[4]
  PIN data_core0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END data_core0[5]
  PIN data_core0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 12.280 75.000 12.880 ;
    END
  END data_core0[6]
  PIN data_core0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END data_core0[7]
  PIN data_core0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END data_core0[8]
  PIN data_core0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 23.160 75.000 23.760 ;
    END
  END data_core0[9]
  PIN is_ready_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END is_ready_core0
  PIN print_hex_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END print_hex_enable
  PIN print_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END print_output[0]
  PIN print_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END print_output[10]
  PIN print_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END print_output[11]
  PIN print_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 71.000 18.770 75.000 ;
    END
  END print_output[12]
  PIN print_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 71.000 27.050 75.000 ;
    END
  END print_output[13]
  PIN print_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END print_output[14]
  PIN print_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 28.600 75.000 29.200 ;
    END
  END print_output[15]
  PIN print_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END print_output[16]
  PIN print_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 39.480 75.000 40.080 ;
    END
  END print_output[17]
  PIN print_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END print_output[18]
  PIN print_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 71.000 39.470 75.000 ;
    END
  END print_output[19]
  PIN print_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END print_output[1]
  PIN print_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END print_output[20]
  PIN print_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 71.000 43.610 75.000 ;
    END
  END print_output[21]
  PIN print_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END print_output[22]
  PIN print_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 71.000 51.890 75.000 ;
    END
  END print_output[23]
  PIN print_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 55.120 75.000 55.720 ;
    END
  END print_output[24]
  PIN print_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END print_output[25]
  PIN print_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 71.000 56.030 75.000 ;
    END
  END print_output[26]
  PIN print_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 71.000 60.170 75.000 ;
    END
  END print_output[27]
  PIN print_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 66.000 75.000 66.600 ;
    END
  END print_output[28]
  PIN print_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 71.000 68.450 75.000 ;
    END
  END print_output[29]
  PIN print_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 6.840 75.000 7.440 ;
    END
  END print_output[2]
  PIN print_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END print_output[30]
  PIN print_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END print_output[31]
  PIN print_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 71.000 10.490 75.000 ;
    END
  END print_output[3]
  PIN print_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END print_output[4]
  PIN print_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 71.000 14.630 75.000 ;
    END
  END print_output[5]
  PIN print_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END print_output[6]
  PIN print_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 17.720 75.000 18.320 ;
    END
  END print_output[7]
  PIN print_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END print_output[8]
  PIN print_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END print_output[9]
  PIN req_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END req_core0
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.380 10.640 16.980 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.700 10.640 38.300 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.020 10.640 59.620 62.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.040 10.640 27.640 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.360 10.640 48.960 62.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 2.465 71.155 62.645 ;
      LAYER met1 ;
        RECT 1.450 2.420 73.070 62.800 ;
      LAYER met2 ;
        RECT 1.480 70.720 1.650 71.925 ;
        RECT 2.490 70.720 5.790 71.925 ;
        RECT 6.630 70.720 9.930 71.925 ;
        RECT 10.770 70.720 14.070 71.925 ;
        RECT 14.910 70.720 18.210 71.925 ;
        RECT 19.050 70.720 22.350 71.925 ;
        RECT 23.190 70.720 26.490 71.925 ;
        RECT 27.330 70.720 30.630 71.925 ;
        RECT 31.470 70.720 34.770 71.925 ;
        RECT 35.610 70.720 38.910 71.925 ;
        RECT 39.750 70.720 43.050 71.925 ;
        RECT 43.890 70.720 47.190 71.925 ;
        RECT 48.030 70.720 51.330 71.925 ;
        RECT 52.170 70.720 55.470 71.925 ;
        RECT 56.310 70.720 59.610 71.925 ;
        RECT 60.450 70.720 63.750 71.925 ;
        RECT 64.590 70.720 67.890 71.925 ;
        RECT 68.730 70.720 72.030 71.925 ;
        RECT 72.870 70.720 73.040 71.925 ;
        RECT 1.480 4.280 73.040 70.720 ;
        RECT 2.030 2.195 4.410 4.280 ;
        RECT 5.250 2.195 8.090 4.280 ;
        RECT 8.930 2.195 11.770 4.280 ;
        RECT 12.610 2.195 15.450 4.280 ;
        RECT 16.290 2.195 18.670 4.280 ;
        RECT 19.510 2.195 22.350 4.280 ;
        RECT 23.190 2.195 26.030 4.280 ;
        RECT 26.870 2.195 29.710 4.280 ;
        RECT 30.550 2.195 32.930 4.280 ;
        RECT 33.770 2.195 36.610 4.280 ;
        RECT 37.450 2.195 40.290 4.280 ;
        RECT 41.130 2.195 43.970 4.280 ;
        RECT 44.810 2.195 47.190 4.280 ;
        RECT 48.030 2.195 50.870 4.280 ;
        RECT 51.710 2.195 54.550 4.280 ;
        RECT 55.390 2.195 58.230 4.280 ;
        RECT 59.070 2.195 61.450 4.280 ;
        RECT 62.290 2.195 65.130 4.280 ;
        RECT 65.970 2.195 68.810 4.280 ;
        RECT 69.650 2.195 72.490 4.280 ;
      LAYER met3 ;
        RECT 4.400 72.440 71.000 72.570 ;
        RECT 4.400 71.720 70.600 72.440 ;
        RECT 4.000 71.040 70.600 71.720 ;
        RECT 4.000 68.360 71.000 71.040 ;
        RECT 4.400 67.000 71.000 68.360 ;
        RECT 4.400 66.960 70.600 67.000 ;
        RECT 4.000 65.600 70.600 66.960 ;
        RECT 4.000 63.600 71.000 65.600 ;
        RECT 4.400 62.200 71.000 63.600 ;
        RECT 4.000 61.560 71.000 62.200 ;
        RECT 4.000 60.160 70.600 61.560 ;
        RECT 4.000 58.840 71.000 60.160 ;
        RECT 4.400 57.440 71.000 58.840 ;
        RECT 4.000 56.120 71.000 57.440 ;
        RECT 4.000 54.720 70.600 56.120 ;
        RECT 4.000 54.080 71.000 54.720 ;
        RECT 4.400 52.680 71.000 54.080 ;
        RECT 4.000 50.680 71.000 52.680 ;
        RECT 4.000 49.320 70.600 50.680 ;
        RECT 4.400 49.280 70.600 49.320 ;
        RECT 4.400 47.920 71.000 49.280 ;
        RECT 4.000 45.240 71.000 47.920 ;
        RECT 4.000 44.560 70.600 45.240 ;
        RECT 4.400 43.840 70.600 44.560 ;
        RECT 4.400 43.160 71.000 43.840 ;
        RECT 4.000 40.480 71.000 43.160 ;
        RECT 4.400 39.080 70.600 40.480 ;
        RECT 4.000 35.720 71.000 39.080 ;
        RECT 4.400 35.040 71.000 35.720 ;
        RECT 4.400 34.320 70.600 35.040 ;
        RECT 4.000 33.640 70.600 34.320 ;
        RECT 4.000 30.960 71.000 33.640 ;
        RECT 4.400 29.600 71.000 30.960 ;
        RECT 4.400 29.560 70.600 29.600 ;
        RECT 4.000 28.200 70.600 29.560 ;
        RECT 4.000 26.200 71.000 28.200 ;
        RECT 4.400 24.800 71.000 26.200 ;
        RECT 4.000 24.160 71.000 24.800 ;
        RECT 4.000 22.760 70.600 24.160 ;
        RECT 4.000 21.440 71.000 22.760 ;
        RECT 4.400 20.040 71.000 21.440 ;
        RECT 4.000 18.720 71.000 20.040 ;
        RECT 4.000 17.320 70.600 18.720 ;
        RECT 4.000 16.680 71.000 17.320 ;
        RECT 4.400 15.280 71.000 16.680 ;
        RECT 4.000 13.280 71.000 15.280 ;
        RECT 4.000 11.920 70.600 13.280 ;
        RECT 4.400 11.880 70.600 11.920 ;
        RECT 4.400 10.520 71.000 11.880 ;
        RECT 4.000 7.840 71.000 10.520 ;
        RECT 4.000 7.160 70.600 7.840 ;
        RECT 4.400 6.440 70.600 7.160 ;
        RECT 4.400 5.760 71.000 6.440 ;
        RECT 4.000 3.080 71.000 5.760 ;
        RECT 4.400 2.215 70.600 3.080 ;
  END
END io_output_arbiter
END LIBRARY

