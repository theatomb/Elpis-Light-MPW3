VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chip_controller
  CLASS BLOCK ;
  FOREIGN chip_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN addr0_to_sram[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END addr0_to_sram[0]
  PIN addr0_to_sram[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 63.280 400.000 63.880 ;
    END
  END addr0_to_sram[10]
  PIN addr0_to_sram[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END addr0_to_sram[11]
  PIN addr0_to_sram[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END addr0_to_sram[12]
  PIN addr0_to_sram[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 78.920 400.000 79.520 ;
    END
  END addr0_to_sram[13]
  PIN addr0_to_sram[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END addr0_to_sram[14]
  PIN addr0_to_sram[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END addr0_to_sram[15]
  PIN addr0_to_sram[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END addr0_to_sram[16]
  PIN addr0_to_sram[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END addr0_to_sram[17]
  PIN addr0_to_sram[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.240 400.000 112.840 ;
    END
  END addr0_to_sram[18]
  PIN addr0_to_sram[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END addr0_to_sram[19]
  PIN addr0_to_sram[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END addr0_to_sram[1]
  PIN addr0_to_sram[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 396.000 16.470 400.000 ;
    END
  END addr0_to_sram[2]
  PIN addr0_to_sram[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 21.120 400.000 21.720 ;
    END
  END addr0_to_sram[3]
  PIN addr0_to_sram[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END addr0_to_sram[4]
  PIN addr0_to_sram[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END addr0_to_sram[5]
  PIN addr0_to_sram[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END addr0_to_sram[6]
  PIN addr0_to_sram[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END addr0_to_sram[7]
  PIN addr0_to_sram[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 396.000 56.490 400.000 ;
    END
  END addr0_to_sram[8]
  PIN addr0_to_sram[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 396.000 68.450 400.000 ;
    END
  END addr0_to_sram[9]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 4.800 400.000 5.400 ;
    END
  END addr_in[0]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END addr_in[10]
  PIN addr_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END addr_in[11]
  PIN addr_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END addr_in[12]
  PIN addr_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 396.000 92.830 400.000 ;
    END
  END addr_in[13]
  PIN addr_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 396.000 97.890 400.000 ;
    END
  END addr_in[14]
  PIN addr_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 89.800 400.000 90.400 ;
    END
  END addr_in[15]
  PIN addr_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END addr_in[16]
  PIN addr_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END addr_in[17]
  PIN addr_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 396.000 125.950 400.000 ;
    END
  END addr_in[18]
  PIN addr_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END addr_in[19]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 12.960 400.000 13.560 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 14.320 400.000 14.920 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 396.000 40.850 400.000 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 41.520 400.000 42.120 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 396.000 50.970 400.000 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 396.000 57.870 400.000 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END addr_in[9]
  PIN addr_to_core_mem[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END addr_to_core_mem[0]
  PIN addr_to_core_mem[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END addr_to_core_mem[10]
  PIN addr_to_core_mem[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END addr_to_core_mem[11]
  PIN addr_to_core_mem[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END addr_to_core_mem[12]
  PIN addr_to_core_mem[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 80.960 400.000 81.560 ;
    END
  END addr_to_core_mem[13]
  PIN addr_to_core_mem[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 82.320 400.000 82.920 ;
    END
  END addr_to_core_mem[14]
  PIN addr_to_core_mem[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 396.000 104.790 400.000 ;
    END
  END addr_to_core_mem[15]
  PIN addr_to_core_mem[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 396.000 112.150 400.000 ;
    END
  END addr_to_core_mem[16]
  PIN addr_to_core_mem[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END addr_to_core_mem[17]
  PIN addr_to_core_mem[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END addr_to_core_mem[18]
  PIN addr_to_core_mem[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 396.000 131.010 400.000 ;
    END
  END addr_to_core_mem[19]
  PIN addr_to_core_mem[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END addr_to_core_mem[1]
  PIN addr_to_core_mem[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END addr_to_core_mem[2]
  PIN addr_to_core_mem[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 396.000 28.430 400.000 ;
    END
  END addr_to_core_mem[3]
  PIN addr_to_core_mem[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 396.000 35.330 400.000 ;
    END
  END addr_to_core_mem[4]
  PIN addr_to_core_mem[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END addr_to_core_mem[5]
  PIN addr_to_core_mem[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 42.880 400.000 43.480 ;
    END
  END addr_to_core_mem[6]
  PIN addr_to_core_mem[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 49.000 400.000 49.600 ;
    END
  END addr_to_core_mem[7]
  PIN addr_to_core_mem[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END addr_to_core_mem[8]
  PIN addr_to_core_mem[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END addr_to_core_mem[9]
  PIN clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END clk
  PIN core0_data_print[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 6.840 400.000 7.440 ;
    END
  END core0_data_print[0]
  PIN core0_data_print[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 64.640 400.000 65.240 ;
    END
  END core0_data_print[10]
  PIN core0_data_print[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END core0_data_print[11]
  PIN core0_data_print[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END core0_data_print[12]
  PIN core0_data_print[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 396.000 94.670 400.000 ;
    END
  END core0_data_print[13]
  PIN core0_data_print[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END core0_data_print[14]
  PIN core0_data_print[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END core0_data_print[15]
  PIN core0_data_print[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END core0_data_print[16]
  PIN core0_data_print[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 396.000 119.050 400.000 ;
    END
  END core0_data_print[17]
  PIN core0_data_print[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 113.600 400.000 114.200 ;
    END
  END core0_data_print[18]
  PIN core0_data_print[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 396.000 132.850 400.000 ;
    END
  END core0_data_print[19]
  PIN core0_data_print[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END core0_data_print[1]
  PIN core0_data_print[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END core0_data_print[20]
  PIN core0_data_print[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END core0_data_print[21]
  PIN core0_data_print[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END core0_data_print[22]
  PIN core0_data_print[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 136.040 400.000 136.640 ;
    END
  END core0_data_print[23]
  PIN core0_data_print[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END core0_data_print[24]
  PIN core0_data_print[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END core0_data_print[25]
  PIN core0_data_print[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END core0_data_print[26]
  PIN core0_data_print[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END core0_data_print[27]
  PIN core0_data_print[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 396.000 183.450 400.000 ;
    END
  END core0_data_print[28]
  PIN core0_data_print[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 163.920 400.000 164.520 ;
    END
  END core0_data_print[29]
  PIN core0_data_print[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 16.360 400.000 16.960 ;
    END
  END core0_data_print[2]
  PIN core0_data_print[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 172.080 400.000 172.680 ;
    END
  END core0_data_print[30]
  PIN core0_data_print[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END core0_data_print[31]
  PIN core0_data_print[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END core0_data_print[3]
  PIN core0_data_print[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 27.240 400.000 27.840 ;
    END
  END core0_data_print[4]
  PIN core0_data_print[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 33.360 400.000 33.960 ;
    END
  END core0_data_print[5]
  PIN core0_data_print[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END core0_data_print[6]
  PIN core0_data_print[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END core0_data_print[7]
  PIN core0_data_print[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 396.000 59.710 400.000 ;
    END
  END core0_data_print[8]
  PIN core0_data_print[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 396.000 70.290 400.000 ;
    END
  END core0_data_print[9]
  PIN csb0_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 2.080 400.000 2.680 ;
    END
  END csb0_to_sram
  PIN data_out_to_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END data_out_to_core[0]
  PIN data_out_to_core[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 396.000 75.350 400.000 ;
    END
  END data_out_to_core[10]
  PIN data_out_to_core[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END data_out_to_core[11]
  PIN data_out_to_core[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 74.160 400.000 74.760 ;
    END
  END data_out_to_core[12]
  PIN data_out_to_core[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END data_out_to_core[13]
  PIN data_out_to_core[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 396.000 99.730 400.000 ;
    END
  END data_out_to_core[14]
  PIN data_out_to_core[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 396.000 106.630 400.000 ;
    END
  END data_out_to_core[15]
  PIN data_out_to_core[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 99.320 400.000 99.920 ;
    END
  END data_out_to_core[16]
  PIN data_out_to_core[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 106.120 400.000 106.720 ;
    END
  END data_out_to_core[17]
  PIN data_out_to_core[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 114.960 400.000 115.560 ;
    END
  END data_out_to_core[18]
  PIN data_out_to_core[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END data_out_to_core[19]
  PIN data_out_to_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END data_out_to_core[1]
  PIN data_out_to_core[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END data_out_to_core[20]
  PIN data_out_to_core[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 396.000 146.650 400.000 ;
    END
  END data_out_to_core[21]
  PIN data_out_to_core[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 396.000 153.550 400.000 ;
    END
  END data_out_to_core[22]
  PIN data_out_to_core[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 396.000 160.910 400.000 ;
    END
  END data_out_to_core[23]
  PIN data_out_to_core[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 396.000 167.810 400.000 ;
    END
  END data_out_to_core[24]
  PIN data_out_to_core[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 396.000 171.030 400.000 ;
    END
  END data_out_to_core[25]
  PIN data_out_to_core[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END data_out_to_core[26]
  PIN data_out_to_core[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END data_out_to_core[27]
  PIN data_out_to_core[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END data_out_to_core[28]
  PIN data_out_to_core[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 165.960 400.000 166.560 ;
    END
  END data_out_to_core[29]
  PIN data_out_to_core[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 396.000 17.850 400.000 ;
    END
  END data_out_to_core[2]
  PIN data_out_to_core[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END data_out_to_core[30]
  PIN data_out_to_core[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 178.200 400.000 178.800 ;
    END
  END data_out_to_core[31]
  PIN data_out_to_core[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 22.480 400.000 23.080 ;
    END
  END data_out_to_core[3]
  PIN data_out_to_core[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END data_out_to_core[4]
  PIN data_out_to_core[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END data_out_to_core[5]
  PIN data_out_to_core[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 44.240 400.000 44.840 ;
    END
  END data_out_to_core[6]
  PIN data_out_to_core[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END data_out_to_core[7]
  PIN data_out_to_core[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END data_out_to_core[8]
  PIN data_out_to_core[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END data_out_to_core[9]
  PIN data_to_core_mem[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 396.000 0.830 400.000 ;
    END
  END data_to_core_mem[0]
  PIN data_to_core_mem[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 66.680 400.000 67.280 ;
    END
  END data_to_core_mem[10]
  PIN data_to_core_mem[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 396.000 82.250 400.000 ;
    END
  END data_to_core_mem[11]
  PIN data_to_core_mem[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 396.000 85.930 400.000 ;
    END
  END data_to_core_mem[12]
  PIN data_to_core_mem[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END data_to_core_mem[13]
  PIN data_to_core_mem[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 83.680 400.000 84.280 ;
    END
  END data_to_core_mem[14]
  PIN data_to_core_mem[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 91.840 400.000 92.440 ;
    END
  END data_to_core_mem[15]
  PIN data_to_core_mem[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 396.000 113.530 400.000 ;
    END
  END data_to_core_mem[16]
  PIN data_to_core_mem[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 107.480 400.000 108.080 ;
    END
  END data_to_core_mem[17]
  PIN data_to_core_mem[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END data_to_core_mem[18]
  PIN data_to_core_mem[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 118.360 400.000 118.960 ;
    END
  END data_to_core_mem[19]
  PIN data_to_core_mem[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END data_to_core_mem[1]
  PIN data_to_core_mem[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 124.480 400.000 125.080 ;
    END
  END data_to_core_mem[20]
  PIN data_to_core_mem[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 396.000 148.490 400.000 ;
    END
  END data_to_core_mem[21]
  PIN data_to_core_mem[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END data_to_core_mem[22]
  PIN data_to_core_mem[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 137.400 400.000 138.000 ;
    END
  END data_to_core_mem[23]
  PIN data_to_core_mem[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 143.520 400.000 144.120 ;
    END
  END data_to_core_mem[24]
  PIN data_to_core_mem[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END data_to_core_mem[25]
  PIN data_to_core_mem[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 153.040 400.000 153.640 ;
    END
  END data_to_core_mem[26]
  PIN data_to_core_mem[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END data_to_core_mem[27]
  PIN data_to_core_mem[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 396.000 184.830 400.000 ;
    END
  END data_to_core_mem[28]
  PIN data_to_core_mem[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END data_to_core_mem[29]
  PIN data_to_core_mem[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 17.720 400.000 18.320 ;
    END
  END data_to_core_mem[2]
  PIN data_to_core_mem[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END data_to_core_mem[30]
  PIN data_to_core_mem[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END data_to_core_mem[31]
  PIN data_to_core_mem[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 396.000 30.270 400.000 ;
    END
  END data_to_core_mem[3]
  PIN data_to_core_mem[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 396.000 37.170 400.000 ;
    END
  END data_to_core_mem[4]
  PIN data_to_core_mem[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 396.000 42.230 400.000 ;
    END
  END data_to_core_mem[5]
  PIN data_to_core_mem[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END data_to_core_mem[6]
  PIN data_to_core_mem[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 51.040 400.000 51.640 ;
    END
  END data_to_core_mem[7]
  PIN data_to_core_mem[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 53.760 400.000 54.360 ;
    END
  END data_to_core_mem[8]
  PIN data_to_core_mem[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END data_to_core_mem[9]
  PIN din0_to_sram[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END din0_to_sram[0]
  PIN din0_to_sram[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 396.000 77.190 400.000 ;
    END
  END din0_to_sram[10]
  PIN din0_to_sram[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END din0_to_sram[11]
  PIN din0_to_sram[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 396.000 87.770 400.000 ;
    END
  END din0_to_sram[12]
  PIN din0_to_sram[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END din0_to_sram[13]
  PIN din0_to_sram[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 85.720 400.000 86.320 ;
    END
  END din0_to_sram[14]
  PIN din0_to_sram[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 396.000 108.470 400.000 ;
    END
  END din0_to_sram[15]
  PIN din0_to_sram[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END din0_to_sram[16]
  PIN din0_to_sram[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END din0_to_sram[17]
  PIN din0_to_sram[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END din0_to_sram[18]
  PIN din0_to_sram[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 119.720 400.000 120.320 ;
    END
  END din0_to_sram[19]
  PIN din0_to_sram[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END din0_to_sram[1]
  PIN din0_to_sram[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END din0_to_sram[20]
  PIN din0_to_sram[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.240 400.000 129.840 ;
    END
  END din0_to_sram[21]
  PIN din0_to_sram[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END din0_to_sram[22]
  PIN din0_to_sram[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END din0_to_sram[23]
  PIN din0_to_sram[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END din0_to_sram[24]
  PIN din0_to_sram[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 396.000 172.870 400.000 ;
    END
  END din0_to_sram[25]
  PIN din0_to_sram[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END din0_to_sram[26]
  PIN din0_to_sram[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 156.440 400.000 157.040 ;
    END
  END din0_to_sram[27]
  PIN din0_to_sram[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END din0_to_sram[28]
  PIN din0_to_sram[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 167.320 400.000 167.920 ;
    END
  END din0_to_sram[29]
  PIN din0_to_sram[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 396.000 19.690 400.000 ;
    END
  END din0_to_sram[2]
  PIN din0_to_sram[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END din0_to_sram[30]
  PIN din0_to_sram[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 179.560 400.000 180.160 ;
    END
  END din0_to_sram[31]
  PIN din0_to_sram[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 23.840 400.000 24.440 ;
    END
  END din0_to_sram[3]
  PIN din0_to_sram[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 396.000 39.010 400.000 ;
    END
  END din0_to_sram[4]
  PIN din0_to_sram[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END din0_to_sram[5]
  PIN din0_to_sram[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END din0_to_sram[6]
  PIN din0_to_sram[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 52.400 400.000 53.000 ;
    END
  END din0_to_sram[7]
  PIN din0_to_sram[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END din0_to_sram[8]
  PIN din0_to_sram[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 57.160 400.000 57.760 ;
    END
  END din0_to_sram[9]
  PIN dout0_to_sram[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 8.200 400.000 8.800 ;
    END
  END dout0_to_sram[0]
  PIN dout0_to_sram[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 396.000 79.030 400.000 ;
    END
  END dout0_to_sram[10]
  PIN dout0_to_sram[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 71.440 400.000 72.040 ;
    END
  END dout0_to_sram[11]
  PIN dout0_to_sram[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 76.200 400.000 76.800 ;
    END
  END dout0_to_sram[12]
  PIN dout0_to_sram[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END dout0_to_sram[13]
  PIN dout0_to_sram[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 87.080 400.000 87.680 ;
    END
  END dout0_to_sram[14]
  PIN dout0_to_sram[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 93.200 400.000 93.800 ;
    END
  END dout0_to_sram[15]
  PIN dout0_to_sram[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 101.360 400.000 101.960 ;
    END
  END dout0_to_sram[16]
  PIN dout0_to_sram[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 396.000 120.890 400.000 ;
    END
  END dout0_to_sram[17]
  PIN dout0_to_sram[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END dout0_to_sram[18]
  PIN dout0_to_sram[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 396.000 134.690 400.000 ;
    END
  END dout0_to_sram[19]
  PIN dout0_to_sram[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 396.000 9.110 400.000 ;
    END
  END dout0_to_sram[1]
  PIN dout0_to_sram[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 396.000 139.750 400.000 ;
    END
  END dout0_to_sram[20]
  PIN dout0_to_sram[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END dout0_to_sram[21]
  PIN dout0_to_sram[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END dout0_to_sram[22]
  PIN dout0_to_sram[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 396.000 162.290 400.000 ;
    END
  END dout0_to_sram[23]
  PIN dout0_to_sram[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END dout0_to_sram[24]
  PIN dout0_to_sram[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END dout0_to_sram[25]
  PIN dout0_to_sram[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END dout0_to_sram[26]
  PIN dout0_to_sram[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END dout0_to_sram[27]
  PIN dout0_to_sram[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 396.000 186.670 400.000 ;
    END
  END dout0_to_sram[28]
  PIN dout0_to_sram[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END dout0_to_sram[29]
  PIN dout0_to_sram[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 19.080 400.000 19.680 ;
    END
  END dout0_to_sram[2]
  PIN dout0_to_sram[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 396.000 195.410 400.000 ;
    END
  END dout0_to_sram[30]
  PIN dout0_to_sram[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 181.600 400.000 182.200 ;
    END
  END dout0_to_sram[31]
  PIN dout0_to_sram[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END dout0_to_sram[3]
  PIN dout0_to_sram[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END dout0_to_sram[4]
  PIN dout0_to_sram[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 34.720 400.000 35.320 ;
    END
  END dout0_to_sram[5]
  PIN dout0_to_sram[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 396.000 45.910 400.000 ;
    END
  END dout0_to_sram[6]
  PIN dout0_to_sram[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END dout0_to_sram[7]
  PIN dout0_to_sram[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END dout0_to_sram[8]
  PIN dout0_to_sram[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 58.520 400.000 59.120 ;
    END
  END dout0_to_sram[9]
  PIN is_loading_memory_into_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END is_loading_memory_into_core
  PIN is_ready_dataout_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END is_ready_dataout_core0
  PIN is_ready_print_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END is_ready_print_core0
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 9.560 400.000 10.160 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 396.000 348.590 400.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 348.200 400.000 348.800 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 396.000 353.650 400.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.720 400.000 358.320 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 396.000 80.870 400.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 396.000 364.230 400.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.520 4.000 348.120 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 396.000 369.290 400.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 378.120 400.000 378.720 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 396.000 378.030 400.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 396.000 379.870 400.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 396.000 390.450 400.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 387.640 400.000 388.240 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 392.400 400.000 393.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 77.560 400.000 78.160 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 94.560 400.000 95.160 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 102.720 400.000 103.320 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 396.000 122.270 400.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 396.000 127.790 400.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 396.000 10.950 400.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 396.000 155.390 400.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 138.760 400.000 139.360 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 396.000 169.190 400.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 148.280 400.000 148.880 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 396.000 176.550 400.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 168.680 400.000 169.280 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 396.000 197.250 400.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 191.120 400.000 191.720 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 195.880 400.000 196.480 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 396.000 211.050 400.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 396.000 214.730 400.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 202.000 400.000 202.600 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.720 400.000 205.320 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 208.120 400.000 208.720 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 396.000 228.530 400.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 219.000 400.000 219.600 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 396.000 240.950 400.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 234.640 400.000 235.240 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 396.000 252.910 400.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 236.680 400.000 237.280 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 396.000 261.650 400.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 396.000 264.870 400.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.920 400.000 249.520 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 396.000 277.290 400.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 396.000 284.190 400.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 264.560 400.000 265.160 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 269.320 400.000 269.920 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 396.000 291.090 400.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 280.880 400.000 281.480 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 396.000 294.770 400.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 288.360 400.000 288.960 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 396.000 52.810 400.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 296.520 400.000 297.120 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 396.000 312.250 400.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 307.400 400.000 308.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 396.000 315.470 400.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 396.000 319.150 400.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 396.000 61.550 400.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 319.640 400.000 320.240 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 326.440 400.000 327.040 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 332.560 400.000 333.160 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 396.000 339.850 400.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 59.880 400.000 60.480 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 396.000 2.210 400.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 343.440 400.000 344.040 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 346.840 400.000 347.440 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 349.560 400.000 350.160 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 352.960 400.000 353.560 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 354.320 400.000 354.920 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 396.000 359.170 400.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 362.480 400.000 363.080 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 396.000 366.070 400.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 370.640 400.000 371.240 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 376.760 400.000 377.360 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 396.000 374.810 400.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 379.480 400.000 380.080 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 381.520 400.000 382.120 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 396.000 381.710 400.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 396.000 384.930 400.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 396.000 392.290 400.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 395.800 400.000 396.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 396.000 89.150 400.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 396.000 96.510 400.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 96.600 400.000 97.200 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 117.000 400.000 117.600 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 396.000 150.330 400.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 396.000 157.230 400.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 144.880 400.000 145.480 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 154.400 400.000 155.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 157.800 400.000 158.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 396.000 188.510 400.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 396.000 192.190 400.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 396.000 21.530 400.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 186.360 400.000 186.960 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 396.000 207.830 400.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 396.000 216.570 400.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 25.880 400.000 26.480 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 203.360 400.000 203.960 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 209.480 400.000 210.080 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 212.880 400.000 213.480 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.040 400.000 221.640 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 396.000 233.590 400.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 396.000 237.270 400.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 396.000 249.230 400.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 396.000 254.750 400.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 239.400 400.000 240.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 241.440 400.000 242.040 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 246.200 400.000 246.800 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 396.000 270.390 400.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 396.000 273.610 400.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 396.000 286.030 400.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 266.600 400.000 267.200 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 46.280 400.000 46.880 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 277.480 400.000 278.080 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 282.240 400.000 282.840 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 396.000 296.610 400.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 396.000 299.830 400.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 293.120 400.000 293.720 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 396.000 303.510 400.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 297.880 400.000 298.480 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 396.000 308.570 400.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 310.800 400.000 311.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 314.880 400.000 315.480 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 396.000 63.390 400.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 396.000 324.210 400.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 324.400 400.000 325.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 396.000 331.110 400.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.920 400.000 334.520 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 335.960 400.000 336.560 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 396.000 334.790 400.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 340.720 400.000 341.320 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 61.920 400.000 62.520 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 396.000 4.050 400.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 344.800 400.000 345.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 396.000 350.430 400.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 396.000 355.490 400.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 361.120 400.000 361.720 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 363.840 400.000 364.440 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.040 400.000 68.640 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 373.360 400.000 373.960 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 396.000 383.550 400.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 389.000 400.000 389.600 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 396.000 395.510 400.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 396.000 115.370 400.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 108.840 400.000 109.440 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 121.760 400.000 122.360 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 396.000 12.790 400.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 126.520 400.000 127.120 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 132.640 400.000 133.240 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 140.800 400.000 141.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 149.640 400.000 150.240 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.160 400.000 159.760 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 173.440 400.000 174.040 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 182.960 400.000 183.560 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 187.720 400.000 188.320 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 396.000 200.930 400.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 396.000 204.150 400.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 396.000 209.210 400.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.240 400.000 197.840 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 396.000 217.950 400.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 396.000 223.470 400.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.240 400.000 214.840 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.280 400.000 216.880 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 396.000 232.210 400.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 396.000 235.430 400.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 396.000 239.110 400.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 396.000 242.330 400.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 28.600 400.000 29.200 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 396.000 244.170 400.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 231.920 400.000 232.520 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 396.000 256.590 400.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 396.000 257.970 400.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 396.000 263.490 400.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 242.800 400.000 243.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 36.760 400.000 37.360 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 396.000 266.710 400.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 255.720 400.000 256.320 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 396.000 279.130 400.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 259.800 400.000 260.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 263.200 400.000 263.800 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 271.360 400.000 271.960 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 274.080 400.000 274.680 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 276.120 400.000 276.720 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 283.600 400.000 284.200 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 289.720 400.000 290.320 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 396.000 304.890 400.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 302.640 400.000 303.240 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 396.000 313.630 400.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 312.160 400.000 312.760 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 396.000 320.990 400.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 396.000 326.050 400.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 327.800 400.000 328.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 329.160 400.000 329.760 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 338.680 400.000 339.280 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 396.000 338.010 400.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 396.000 341.690 400.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END la_oenb[9]
  PIN rd_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END rd_data_out[0]
  PIN rd_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END rd_data_out[100]
  PIN rd_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END rd_data_out[101]
  PIN rd_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END rd_data_out[102]
  PIN rd_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END rd_data_out[103]
  PIN rd_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 396.000 357.330 400.000 ;
    END
  END rd_data_out[104]
  PIN rd_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END rd_data_out[105]
  PIN rd_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 356.360 400.000 356.960 ;
    END
  END rd_data_out[106]
  PIN rd_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END rd_data_out[107]
  PIN rd_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END rd_data_out[108]
  PIN rd_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 396.000 362.390 400.000 ;
    END
  END rd_data_out[109]
  PIN rd_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END rd_data_out[10]
  PIN rd_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 367.240 400.000 367.840 ;
    END
  END rd_data_out[110]
  PIN rd_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END rd_data_out[111]
  PIN rd_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END rd_data_out[112]
  PIN rd_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 396.000 367.910 400.000 ;
    END
  END rd_data_out[113]
  PIN rd_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 396.000 371.130 400.000 ;
    END
  END rd_data_out[114]
  PIN rd_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 396.000 372.970 400.000 ;
    END
  END rd_data_out[115]
  PIN rd_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END rd_data_out[116]
  PIN rd_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 396.000 376.650 400.000 ;
    END
  END rd_data_out[117]
  PIN rd_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END rd_data_out[118]
  PIN rd_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END rd_data_out[119]
  PIN rd_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END rd_data_out[11]
  PIN rd_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END rd_data_out[120]
  PIN rd_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 382.880 400.000 383.480 ;
    END
  END rd_data_out[121]
  PIN rd_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 396.000 386.770 400.000 ;
    END
  END rd_data_out[122]
  PIN rd_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END rd_data_out[123]
  PIN rd_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 396.000 393.670 400.000 ;
    END
  END rd_data_out[124]
  PIN rd_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 396.000 397.350 400.000 ;
    END
  END rd_data_out[125]
  PIN rd_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 397.160 400.000 397.760 ;
    END
  END rd_data_out[126]
  PIN rd_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END rd_data_out[127]
  PIN rd_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 396.000 90.990 400.000 ;
    END
  END rd_data_out[12]
  PIN rd_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END rd_data_out[13]
  PIN rd_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 88.440 400.000 89.040 ;
    END
  END rd_data_out[14]
  PIN rd_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 396.000 110.310 400.000 ;
    END
  END rd_data_out[15]
  PIN rd_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 104.080 400.000 104.680 ;
    END
  END rd_data_out[16]
  PIN rd_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 110.880 400.000 111.480 ;
    END
  END rd_data_out[17]
  PIN rd_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END rd_data_out[18]
  PIN rd_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 396.000 136.530 400.000 ;
    END
  END rd_data_out[19]
  PIN rd_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END rd_data_out[1]
  PIN rd_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 396.000 141.590 400.000 ;
    END
  END rd_data_out[20]
  PIN rd_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END rd_data_out[21]
  PIN rd_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END rd_data_out[22]
  PIN rd_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 396.000 164.130 400.000 ;
    END
  END rd_data_out[23]
  PIN rd_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END rd_data_out[24]
  PIN rd_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END rd_data_out[25]
  PIN rd_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 396.000 177.930 400.000 ;
    END
  END rd_data_out[26]
  PIN rd_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 396.000 181.610 400.000 ;
    END
  END rd_data_out[27]
  PIN rd_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END rd_data_out[28]
  PIN rd_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 396.000 193.570 400.000 ;
    END
  END rd_data_out[29]
  PIN rd_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END rd_data_out[2]
  PIN rd_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END rd_data_out[30]
  PIN rd_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END rd_data_out[31]
  PIN rd_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 189.080 400.000 189.680 ;
    END
  END rd_data_out[32]
  PIN rd_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 396.000 202.310 400.000 ;
    END
  END rd_data_out[33]
  PIN rd_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END rd_data_out[34]
  PIN rd_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 396.000 205.990 400.000 ;
    END
  END rd_data_out[35]
  PIN rd_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END rd_data_out[36]
  PIN rd_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 396.000 212.890 400.000 ;
    END
  END rd_data_out[37]
  PIN rd_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END rd_data_out[38]
  PIN rd_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 200.640 400.000 201.240 ;
    END
  END rd_data_out[39]
  PIN rd_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END rd_data_out[3]
  PIN rd_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END rd_data_out[40]
  PIN rd_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 396.000 221.630 400.000 ;
    END
  END rd_data_out[41]
  PIN rd_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END rd_data_out[42]
  PIN rd_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 396.000 224.850 400.000 ;
    END
  END rd_data_out[43]
  PIN rd_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END rd_data_out[44]
  PIN rd_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 217.640 400.000 218.240 ;
    END
  END rd_data_out[45]
  PIN rd_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 222.400 400.000 223.000 ;
    END
  END rd_data_out[46]
  PIN rd_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 223.760 400.000 224.360 ;
    END
  END rd_data_out[47]
  PIN rd_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END rd_data_out[48]
  PIN rd_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END rd_data_out[49]
  PIN rd_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END rd_data_out[4]
  PIN rd_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 228.520 400.000 229.120 ;
    END
  END rd_data_out[50]
  PIN rd_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END rd_data_out[51]
  PIN rd_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 396.000 247.850 400.000 ;
    END
  END rd_data_out[52]
  PIN rd_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END rd_data_out[53]
  PIN rd_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END rd_data_out[54]
  PIN rd_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END rd_data_out[55]
  PIN rd_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END rd_data_out[56]
  PIN rd_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.040 400.000 238.640 ;
    END
  END rd_data_out[57]
  PIN rd_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END rd_data_out[58]
  PIN rd_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 244.160 400.000 244.760 ;
    END
  END rd_data_out[59]
  PIN rd_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 396.000 44.070 400.000 ;
    END
  END rd_data_out[5]
  PIN rd_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 396.000 268.550 400.000 ;
    END
  END rd_data_out[60]
  PIN rd_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 250.960 400.000 251.560 ;
    END
  END rd_data_out[61]
  PIN rd_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 252.320 400.000 252.920 ;
    END
  END rd_data_out[62]
  PIN rd_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 396.000 272.230 400.000 ;
    END
  END rd_data_out[63]
  PIN rd_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 258.440 400.000 259.040 ;
    END
  END rd_data_out[64]
  PIN rd_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 396.000 280.970 400.000 ;
    END
  END rd_data_out[65]
  PIN rd_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END rd_data_out[66]
  PIN rd_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END rd_data_out[67]
  PIN rd_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 267.960 400.000 268.560 ;
    END
  END rd_data_out[68]
  PIN rd_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END rd_data_out[69]
  PIN rd_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 396.000 47.750 400.000 ;
    END
  END rd_data_out[6]
  PIN rd_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END rd_data_out[70]
  PIN rd_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 396.000 289.250 400.000 ;
    END
  END rd_data_out[71]
  PIN rd_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END rd_data_out[72]
  PIN rd_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.840 400.000 279.440 ;
    END
  END rd_data_out[73]
  PIN rd_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 285.640 400.000 286.240 ;
    END
  END rd_data_out[74]
  PIN rd_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END rd_data_out[75]
  PIN rd_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 291.760 400.000 292.360 ;
    END
  END rd_data_out[76]
  PIN rd_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END rd_data_out[77]
  PIN rd_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END rd_data_out[78]
  PIN rd_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 294.480 400.000 295.080 ;
    END
  END rd_data_out[79]
  PIN rd_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 396.000 54.650 400.000 ;
    END
  END rd_data_out[7]
  PIN rd_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 299.240 400.000 299.840 ;
    END
  END rd_data_out[80]
  PIN rd_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 396.000 310.410 400.000 ;
    END
  END rd_data_out[81]
  PIN rd_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 301.280 400.000 301.880 ;
    END
  END rd_data_out[82]
  PIN rd_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 304.000 400.000 304.600 ;
    END
  END rd_data_out[83]
  PIN rd_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END rd_data_out[84]
  PIN rd_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END rd_data_out[85]
  PIN rd_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END rd_data_out[86]
  PIN rd_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 396.000 317.310 400.000 ;
    END
  END rd_data_out[87]
  PIN rd_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 316.920 400.000 317.520 ;
    END
  END rd_data_out[88]
  PIN rd_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 318.280 400.000 318.880 ;
    END
  END rd_data_out[89]
  PIN rd_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END rd_data_out[8]
  PIN rd_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END rd_data_out[90]
  PIN rd_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END rd_data_out[91]
  PIN rd_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 396.000 327.890 400.000 ;
    END
  END rd_data_out[92]
  PIN rd_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 396.000 329.270 400.000 ;
    END
  END rd_data_out[93]
  PIN rd_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END rd_data_out[94]
  PIN rd_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END rd_data_out[95]
  PIN rd_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 396.000 332.950 400.000 ;
    END
  END rd_data_out[96]
  PIN rd_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 396.000 336.630 400.000 ;
    END
  END rd_data_out[97]
  PIN rd_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 342.080 400.000 342.680 ;
    END
  END rd_data_out[98]
  PIN rd_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 396.000 343.530 400.000 ;
    END
  END rd_data_out[99]
  PIN rd_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END rd_data_out[9]
  PIN read_enable_to_Elpis
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END read_enable_to_Elpis
  PIN read_interactive_req_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END read_interactive_req_core0
  PIN read_value_to_Elpis[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 11.600 400.000 12.200 ;
    END
  END read_value_to_Elpis[0]
  PIN read_value_to_Elpis[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END read_value_to_Elpis[10]
  PIN read_value_to_Elpis[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 396.000 84.090 400.000 ;
    END
  END read_value_to_Elpis[11]
  PIN read_value_to_Elpis[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END read_value_to_Elpis[12]
  PIN read_value_to_Elpis[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END read_value_to_Elpis[13]
  PIN read_value_to_Elpis[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END read_value_to_Elpis[14]
  PIN read_value_to_Elpis[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 97.960 400.000 98.560 ;
    END
  END read_value_to_Elpis[15]
  PIN read_value_to_Elpis[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 396.000 117.210 400.000 ;
    END
  END read_value_to_Elpis[16]
  PIN read_value_to_Elpis[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END read_value_to_Elpis[17]
  PIN read_value_to_Elpis[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 396.000 129.170 400.000 ;
    END
  END read_value_to_Elpis[18]
  PIN read_value_to_Elpis[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END read_value_to_Elpis[19]
  PIN read_value_to_Elpis[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 396.000 14.630 400.000 ;
    END
  END read_value_to_Elpis[1]
  PIN read_value_to_Elpis[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 127.880 400.000 128.480 ;
    END
  END read_value_to_Elpis[20]
  PIN read_value_to_Elpis[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 396.000 152.170 400.000 ;
    END
  END read_value_to_Elpis[21]
  PIN read_value_to_Elpis[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 396.000 159.070 400.000 ;
    END
  END read_value_to_Elpis[22]
  PIN read_value_to_Elpis[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.160 400.000 142.760 ;
    END
  END read_value_to_Elpis[23]
  PIN read_value_to_Elpis[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 146.920 400.000 147.520 ;
    END
  END read_value_to_Elpis[24]
  PIN read_value_to_Elpis[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 396.000 174.710 400.000 ;
    END
  END read_value_to_Elpis[25]
  PIN read_value_to_Elpis[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END read_value_to_Elpis[26]
  PIN read_value_to_Elpis[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END read_value_to_Elpis[27]
  PIN read_value_to_Elpis[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 396.000 190.350 400.000 ;
    END
  END read_value_to_Elpis[28]
  PIN read_value_to_Elpis[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END read_value_to_Elpis[29]
  PIN read_value_to_Elpis[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 396.000 23.370 400.000 ;
    END
  END read_value_to_Elpis[2]
  PIN read_value_to_Elpis[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END read_value_to_Elpis[30]
  PIN read_value_to_Elpis[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END read_value_to_Elpis[31]
  PIN read_value_to_Elpis[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 396.000 32.110 400.000 ;
    END
  END read_value_to_Elpis[3]
  PIN read_value_to_Elpis[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END read_value_to_Elpis[4]
  PIN read_value_to_Elpis[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END read_value_to_Elpis[5]
  PIN read_value_to_Elpis[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 47.640 400.000 48.240 ;
    END
  END read_value_to_Elpis[6]
  PIN read_value_to_Elpis[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END read_value_to_Elpis[7]
  PIN read_value_to_Elpis[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 396.000 64.770 400.000 ;
    END
  END read_value_to_Elpis[8]
  PIN read_value_to_Elpis[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 396.000 72.130 400.000 ;
    END
  END read_value_to_Elpis[9]
  PIN ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END ready
  PIN req_out_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END req_out_core0
  PIN requested
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END requested
  PIN reset_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END reset_core
  PIN reset_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END reset_mem_req
  PIN rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END rst
  PIN spare_wen0_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 3.440 400.000 4.040 ;
    END
  END spare_wen0_to_sram
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_rst_i
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 396.000 5.890 400.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 69.400 400.000 70.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 396.000 101.570 400.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 396.000 137.910 400.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 396.000 143.430 400.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 151.680 400.000 152.280 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 396.000 179.770 400.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 161.200 400.000 161.800 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.720 400.000 171.320 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 396.000 24.750 400.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 174.800 400.000 175.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 396.000 199.090 400.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 29.960 400.000 30.560 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 38.120 400.000 38.720 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 396.000 49.130 400.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 55.800 400.000 56.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 396.000 73.510 400.000 ;
    END
  END wbs_dat_o[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END we
  PIN we_to_sram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 0.720 400.000 1.320 ;
    END
  END we_to_sram
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 396.000 7.730 400.000 ;
    END
  END wr_data[0]
  PIN wr_data[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 396.000 346.750 400.000 ;
    END
  END wr_data[100]
  PIN wr_data[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 396.000 352.270 400.000 ;
    END
  END wr_data[101]
  PIN wr_data[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 351.600 400.000 352.200 ;
    END
  END wr_data[102]
  PIN wr_data[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END wr_data[103]
  PIN wr_data[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END wr_data[104]
  PIN wr_data[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END wr_data[105]
  PIN wr_data[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END wr_data[106]
  PIN wr_data[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 359.080 400.000 359.680 ;
    END
  END wr_data[107]
  PIN wr_data[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 396.000 361.010 400.000 ;
    END
  END wr_data[108]
  PIN wr_data[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 365.880 400.000 366.480 ;
    END
  END wr_data[109]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END wr_data[10]
  PIN wr_data[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 368.600 400.000 369.200 ;
    END
  END wr_data[110]
  PIN wr_data[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 372.000 400.000 372.600 ;
    END
  END wr_data[111]
  PIN wr_data[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END wr_data[112]
  PIN wr_data[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END wr_data[113]
  PIN wr_data[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 374.720 400.000 375.320 ;
    END
  END wr_data[114]
  PIN wr_data[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END wr_data[115]
  PIN wr_data[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END wr_data[116]
  PIN wr_data[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END wr_data[117]
  PIN wr_data[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END wr_data[118]
  PIN wr_data[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END wr_data[119]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 72.800 400.000 73.400 ;
    END
  END wr_data[11]
  PIN wr_data[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END wr_data[120]
  PIN wr_data[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 384.240 400.000 384.840 ;
    END
  END wr_data[121]
  PIN wr_data[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 396.000 388.610 400.000 ;
    END
  END wr_data[122]
  PIN wr_data[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 386.280 400.000 386.880 ;
    END
  END wr_data[123]
  PIN wr_data[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 391.040 400.000 391.640 ;
    END
  END wr_data[124]
  PIN wr_data[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 393.760 400.000 394.360 ;
    END
  END wr_data[125]
  PIN wr_data[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 398.520 400.000 399.120 ;
    END
  END wr_data[126]
  PIN wr_data[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 396.000 399.190 400.000 ;
    END
  END wr_data[127]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END wr_data[12]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wr_data[13]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 396.000 103.410 400.000 ;
    END
  END wr_data[14]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END wr_data[15]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wr_data[16]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 396.000 124.110 400.000 ;
    END
  END wr_data[17]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wr_data[18]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.120 400.000 123.720 ;
    END
  END wr_data[19]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END wr_data[1]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 396.000 144.810 400.000 ;
    END
  END wr_data[20]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 131.280 400.000 131.880 ;
    END
  END wr_data[21]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 134.000 400.000 134.600 ;
    END
  END wr_data[22]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 396.000 165.970 400.000 ;
    END
  END wr_data[23]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wr_data[24]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wr_data[25]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END wr_data[26]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END wr_data[27]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 162.560 400.000 163.160 ;
    END
  END wr_data[28]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END wr_data[29]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 396.000 26.590 400.000 ;
    END
  END wr_data[2]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 176.840 400.000 177.440 ;
    END
  END wr_data[30]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 184.320 400.000 184.920 ;
    END
  END wr_data[31]
  PIN wr_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END wr_data[32]
  PIN wr_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wr_data[33]
  PIN wr_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 192.480 400.000 193.080 ;
    END
  END wr_data[34]
  PIN wr_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.840 400.000 194.440 ;
    END
  END wr_data[35]
  PIN wr_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END wr_data[36]
  PIN wr_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END wr_data[37]
  PIN wr_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 198.600 400.000 199.200 ;
    END
  END wr_data[38]
  PIN wr_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END wr_data[39]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 396.000 33.490 400.000 ;
    END
  END wr_data[3]
  PIN wr_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 396.000 219.790 400.000 ;
    END
  END wr_data[40]
  PIN wr_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END wr_data[41]
  PIN wr_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 206.760 400.000 207.360 ;
    END
  END wr_data[42]
  PIN wr_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 211.520 400.000 212.120 ;
    END
  END wr_data[43]
  PIN wr_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 396.000 226.690 400.000 ;
    END
  END wr_data[44]
  PIN wr_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 396.000 230.370 400.000 ;
    END
  END wr_data[45]
  PIN wr_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END wr_data[46]
  PIN wr_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END wr_data[47]
  PIN wr_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 225.800 400.000 226.400 ;
    END
  END wr_data[48]
  PIN wr_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.160 400.000 227.760 ;
    END
  END wr_data[49]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 32.000 400.000 32.600 ;
    END
  END wr_data[4]
  PIN wr_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 229.880 400.000 230.480 ;
    END
  END wr_data[50]
  PIN wr_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 396.000 246.010 400.000 ;
    END
  END wr_data[51]
  PIN wr_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 233.280 400.000 233.880 ;
    END
  END wr_data[52]
  PIN wr_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 396.000 251.070 400.000 ;
    END
  END wr_data[53]
  PIN wr_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END wr_data[54]
  PIN wr_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END wr_data[55]
  PIN wr_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 396.000 259.810 400.000 ;
    END
  END wr_data[56]
  PIN wr_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END wr_data[57]
  PIN wr_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END wr_data[58]
  PIN wr_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END wr_data[59]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 39.480 400.000 40.080 ;
    END
  END wr_data[5]
  PIN wr_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 247.560 400.000 248.160 ;
    END
  END wr_data[60]
  PIN wr_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END wr_data[61]
  PIN wr_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 253.680 400.000 254.280 ;
    END
  END wr_data[62]
  PIN wr_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 257.080 400.000 257.680 ;
    END
  END wr_data[63]
  PIN wr_data[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 396.000 275.450 400.000 ;
    END
  END wr_data[64]
  PIN wr_data[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 396.000 282.350 400.000 ;
    END
  END wr_data[65]
  PIN wr_data[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 261.840 400.000 262.440 ;
    END
  END wr_data[66]
  PIN wr_data[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 396.000 287.870 400.000 ;
    END
  END wr_data[67]
  PIN wr_data[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END wr_data[68]
  PIN wr_data[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 272.720 400.000 273.320 ;
    END
  END wr_data[69]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wr_data[6]
  PIN wr_data[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wr_data[70]
  PIN wr_data[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END wr_data[71]
  PIN wr_data[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END wr_data[72]
  PIN wr_data[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 396.000 292.930 400.000 ;
    END
  END wr_data[73]
  PIN wr_data[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 287.000 400.000 287.600 ;
    END
  END wr_data[74]
  PIN wr_data[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 396.000 297.990 400.000 ;
    END
  END wr_data[75]
  PIN wr_data[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END wr_data[76]
  PIN wr_data[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 396.000 301.670 400.000 ;
    END
  END wr_data[77]
  PIN wr_data[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END wr_data[78]
  PIN wr_data[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END wr_data[79]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END wr_data[7]
  PIN wr_data[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 396.000 306.730 400.000 ;
    END
  END wr_data[80]
  PIN wr_data[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END wr_data[81]
  PIN wr_data[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END wr_data[82]
  PIN wr_data[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.040 400.000 306.640 ;
    END
  END wr_data[83]
  PIN wr_data[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 308.760 400.000 309.360 ;
    END
  END wr_data[84]
  PIN wr_data[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END wr_data[85]
  PIN wr_data[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END wr_data[86]
  PIN wr_data[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 313.520 400.000 314.120 ;
    END
  END wr_data[87]
  PIN wr_data[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END wr_data[88]
  PIN wr_data[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 396.000 322.370 400.000 ;
    END
  END wr_data[89]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 396.000 66.610 400.000 ;
    END
  END wr_data[8]
  PIN wr_data[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.680 400.000 322.280 ;
    END
  END wr_data[90]
  PIN wr_data[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 323.040 400.000 323.640 ;
    END
  END wr_data[91]
  PIN wr_data[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END wr_data[92]
  PIN wr_data[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END wr_data[93]
  PIN wr_data[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 331.200 400.000 331.800 ;
    END
  END wr_data[94]
  PIN wr_data[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END wr_data[95]
  PIN wr_data[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 337.320 400.000 337.920 ;
    END
  END wr_data[96]
  PIN wr_data[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END wr_data[97]
  PIN wr_data[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END wr_data[98]
  PIN wr_data[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 396.000 344.910 400.000 ;
    END
  END wr_data[99]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END wr_data[9]
  OBS
      LAYER li1 ;
        RECT 5.520 5.185 396.835 393.975 ;
      LAYER met1 ;
        RECT 0.530 5.140 399.210 394.020 ;
      LAYER met2 ;
        RECT 1.110 395.720 1.650 399.005 ;
        RECT 2.490 395.720 3.490 399.005 ;
        RECT 4.330 395.720 5.330 399.005 ;
        RECT 6.170 395.720 7.170 399.005 ;
        RECT 8.010 395.720 8.550 399.005 ;
        RECT 9.390 395.720 10.390 399.005 ;
        RECT 11.230 395.720 12.230 399.005 ;
        RECT 13.070 395.720 14.070 399.005 ;
        RECT 14.910 395.720 15.910 399.005 ;
        RECT 16.750 395.720 17.290 399.005 ;
        RECT 18.130 395.720 19.130 399.005 ;
        RECT 19.970 395.720 20.970 399.005 ;
        RECT 21.810 395.720 22.810 399.005 ;
        RECT 23.650 395.720 24.190 399.005 ;
        RECT 25.030 395.720 26.030 399.005 ;
        RECT 26.870 395.720 27.870 399.005 ;
        RECT 28.710 395.720 29.710 399.005 ;
        RECT 30.550 395.720 31.550 399.005 ;
        RECT 32.390 395.720 32.930 399.005 ;
        RECT 33.770 395.720 34.770 399.005 ;
        RECT 35.610 395.720 36.610 399.005 ;
        RECT 37.450 395.720 38.450 399.005 ;
        RECT 39.290 395.720 40.290 399.005 ;
        RECT 41.130 395.720 41.670 399.005 ;
        RECT 42.510 395.720 43.510 399.005 ;
        RECT 44.350 395.720 45.350 399.005 ;
        RECT 46.190 395.720 47.190 399.005 ;
        RECT 48.030 395.720 48.570 399.005 ;
        RECT 49.410 395.720 50.410 399.005 ;
        RECT 51.250 395.720 52.250 399.005 ;
        RECT 53.090 395.720 54.090 399.005 ;
        RECT 54.930 395.720 55.930 399.005 ;
        RECT 56.770 395.720 57.310 399.005 ;
        RECT 58.150 395.720 59.150 399.005 ;
        RECT 59.990 395.720 60.990 399.005 ;
        RECT 61.830 395.720 62.830 399.005 ;
        RECT 63.670 395.720 64.210 399.005 ;
        RECT 65.050 395.720 66.050 399.005 ;
        RECT 66.890 395.720 67.890 399.005 ;
        RECT 68.730 395.720 69.730 399.005 ;
        RECT 70.570 395.720 71.570 399.005 ;
        RECT 72.410 395.720 72.950 399.005 ;
        RECT 73.790 395.720 74.790 399.005 ;
        RECT 75.630 395.720 76.630 399.005 ;
        RECT 77.470 395.720 78.470 399.005 ;
        RECT 79.310 395.720 80.310 399.005 ;
        RECT 81.150 395.720 81.690 399.005 ;
        RECT 82.530 395.720 83.530 399.005 ;
        RECT 84.370 395.720 85.370 399.005 ;
        RECT 86.210 395.720 87.210 399.005 ;
        RECT 88.050 395.720 88.590 399.005 ;
        RECT 89.430 395.720 90.430 399.005 ;
        RECT 91.270 395.720 92.270 399.005 ;
        RECT 93.110 395.720 94.110 399.005 ;
        RECT 94.950 395.720 95.950 399.005 ;
        RECT 96.790 395.720 97.330 399.005 ;
        RECT 98.170 395.720 99.170 399.005 ;
        RECT 100.010 395.720 101.010 399.005 ;
        RECT 101.850 395.720 102.850 399.005 ;
        RECT 103.690 395.720 104.230 399.005 ;
        RECT 105.070 395.720 106.070 399.005 ;
        RECT 106.910 395.720 107.910 399.005 ;
        RECT 108.750 395.720 109.750 399.005 ;
        RECT 110.590 395.720 111.590 399.005 ;
        RECT 112.430 395.720 112.970 399.005 ;
        RECT 113.810 395.720 114.810 399.005 ;
        RECT 115.650 395.720 116.650 399.005 ;
        RECT 117.490 395.720 118.490 399.005 ;
        RECT 119.330 395.720 120.330 399.005 ;
        RECT 121.170 395.720 121.710 399.005 ;
        RECT 122.550 395.720 123.550 399.005 ;
        RECT 124.390 395.720 125.390 399.005 ;
        RECT 126.230 395.720 127.230 399.005 ;
        RECT 128.070 395.720 128.610 399.005 ;
        RECT 129.450 395.720 130.450 399.005 ;
        RECT 131.290 395.720 132.290 399.005 ;
        RECT 133.130 395.720 134.130 399.005 ;
        RECT 134.970 395.720 135.970 399.005 ;
        RECT 136.810 395.720 137.350 399.005 ;
        RECT 138.190 395.720 139.190 399.005 ;
        RECT 140.030 395.720 141.030 399.005 ;
        RECT 141.870 395.720 142.870 399.005 ;
        RECT 143.710 395.720 144.250 399.005 ;
        RECT 145.090 395.720 146.090 399.005 ;
        RECT 146.930 395.720 147.930 399.005 ;
        RECT 148.770 395.720 149.770 399.005 ;
        RECT 150.610 395.720 151.610 399.005 ;
        RECT 152.450 395.720 152.990 399.005 ;
        RECT 153.830 395.720 154.830 399.005 ;
        RECT 155.670 395.720 156.670 399.005 ;
        RECT 157.510 395.720 158.510 399.005 ;
        RECT 159.350 395.720 160.350 399.005 ;
        RECT 161.190 395.720 161.730 399.005 ;
        RECT 162.570 395.720 163.570 399.005 ;
        RECT 164.410 395.720 165.410 399.005 ;
        RECT 166.250 395.720 167.250 399.005 ;
        RECT 168.090 395.720 168.630 399.005 ;
        RECT 169.470 395.720 170.470 399.005 ;
        RECT 171.310 395.720 172.310 399.005 ;
        RECT 173.150 395.720 174.150 399.005 ;
        RECT 174.990 395.720 175.990 399.005 ;
        RECT 176.830 395.720 177.370 399.005 ;
        RECT 178.210 395.720 179.210 399.005 ;
        RECT 180.050 395.720 181.050 399.005 ;
        RECT 181.890 395.720 182.890 399.005 ;
        RECT 183.730 395.720 184.270 399.005 ;
        RECT 185.110 395.720 186.110 399.005 ;
        RECT 186.950 395.720 187.950 399.005 ;
        RECT 188.790 395.720 189.790 399.005 ;
        RECT 190.630 395.720 191.630 399.005 ;
        RECT 192.470 395.720 193.010 399.005 ;
        RECT 193.850 395.720 194.850 399.005 ;
        RECT 195.690 395.720 196.690 399.005 ;
        RECT 197.530 395.720 198.530 399.005 ;
        RECT 199.370 395.720 200.370 399.005 ;
        RECT 201.210 395.720 201.750 399.005 ;
        RECT 202.590 395.720 203.590 399.005 ;
        RECT 204.430 395.720 205.430 399.005 ;
        RECT 206.270 395.720 207.270 399.005 ;
        RECT 208.110 395.720 208.650 399.005 ;
        RECT 209.490 395.720 210.490 399.005 ;
        RECT 211.330 395.720 212.330 399.005 ;
        RECT 213.170 395.720 214.170 399.005 ;
        RECT 215.010 395.720 216.010 399.005 ;
        RECT 216.850 395.720 217.390 399.005 ;
        RECT 218.230 395.720 219.230 399.005 ;
        RECT 220.070 395.720 221.070 399.005 ;
        RECT 221.910 395.720 222.910 399.005 ;
        RECT 223.750 395.720 224.290 399.005 ;
        RECT 225.130 395.720 226.130 399.005 ;
        RECT 226.970 395.720 227.970 399.005 ;
        RECT 228.810 395.720 229.810 399.005 ;
        RECT 230.650 395.720 231.650 399.005 ;
        RECT 232.490 395.720 233.030 399.005 ;
        RECT 233.870 395.720 234.870 399.005 ;
        RECT 235.710 395.720 236.710 399.005 ;
        RECT 237.550 395.720 238.550 399.005 ;
        RECT 239.390 395.720 240.390 399.005 ;
        RECT 241.230 395.720 241.770 399.005 ;
        RECT 242.610 395.720 243.610 399.005 ;
        RECT 244.450 395.720 245.450 399.005 ;
        RECT 246.290 395.720 247.290 399.005 ;
        RECT 248.130 395.720 248.670 399.005 ;
        RECT 249.510 395.720 250.510 399.005 ;
        RECT 251.350 395.720 252.350 399.005 ;
        RECT 253.190 395.720 254.190 399.005 ;
        RECT 255.030 395.720 256.030 399.005 ;
        RECT 256.870 395.720 257.410 399.005 ;
        RECT 258.250 395.720 259.250 399.005 ;
        RECT 260.090 395.720 261.090 399.005 ;
        RECT 261.930 395.720 262.930 399.005 ;
        RECT 263.770 395.720 264.310 399.005 ;
        RECT 265.150 395.720 266.150 399.005 ;
        RECT 266.990 395.720 267.990 399.005 ;
        RECT 268.830 395.720 269.830 399.005 ;
        RECT 270.670 395.720 271.670 399.005 ;
        RECT 272.510 395.720 273.050 399.005 ;
        RECT 273.890 395.720 274.890 399.005 ;
        RECT 275.730 395.720 276.730 399.005 ;
        RECT 277.570 395.720 278.570 399.005 ;
        RECT 279.410 395.720 280.410 399.005 ;
        RECT 281.250 395.720 281.790 399.005 ;
        RECT 282.630 395.720 283.630 399.005 ;
        RECT 284.470 395.720 285.470 399.005 ;
        RECT 286.310 395.720 287.310 399.005 ;
        RECT 288.150 395.720 288.690 399.005 ;
        RECT 289.530 395.720 290.530 399.005 ;
        RECT 291.370 395.720 292.370 399.005 ;
        RECT 293.210 395.720 294.210 399.005 ;
        RECT 295.050 395.720 296.050 399.005 ;
        RECT 296.890 395.720 297.430 399.005 ;
        RECT 298.270 395.720 299.270 399.005 ;
        RECT 300.110 395.720 301.110 399.005 ;
        RECT 301.950 395.720 302.950 399.005 ;
        RECT 303.790 395.720 304.330 399.005 ;
        RECT 305.170 395.720 306.170 399.005 ;
        RECT 307.010 395.720 308.010 399.005 ;
        RECT 308.850 395.720 309.850 399.005 ;
        RECT 310.690 395.720 311.690 399.005 ;
        RECT 312.530 395.720 313.070 399.005 ;
        RECT 313.910 395.720 314.910 399.005 ;
        RECT 315.750 395.720 316.750 399.005 ;
        RECT 317.590 395.720 318.590 399.005 ;
        RECT 319.430 395.720 320.430 399.005 ;
        RECT 321.270 395.720 321.810 399.005 ;
        RECT 322.650 395.720 323.650 399.005 ;
        RECT 324.490 395.720 325.490 399.005 ;
        RECT 326.330 395.720 327.330 399.005 ;
        RECT 328.170 395.720 328.710 399.005 ;
        RECT 329.550 395.720 330.550 399.005 ;
        RECT 331.390 395.720 332.390 399.005 ;
        RECT 333.230 395.720 334.230 399.005 ;
        RECT 335.070 395.720 336.070 399.005 ;
        RECT 336.910 395.720 337.450 399.005 ;
        RECT 338.290 395.720 339.290 399.005 ;
        RECT 340.130 395.720 341.130 399.005 ;
        RECT 341.970 395.720 342.970 399.005 ;
        RECT 343.810 395.720 344.350 399.005 ;
        RECT 345.190 395.720 346.190 399.005 ;
        RECT 347.030 395.720 348.030 399.005 ;
        RECT 348.870 395.720 349.870 399.005 ;
        RECT 350.710 395.720 351.710 399.005 ;
        RECT 352.550 395.720 353.090 399.005 ;
        RECT 353.930 395.720 354.930 399.005 ;
        RECT 355.770 395.720 356.770 399.005 ;
        RECT 357.610 395.720 358.610 399.005 ;
        RECT 359.450 395.720 360.450 399.005 ;
        RECT 361.290 395.720 361.830 399.005 ;
        RECT 362.670 395.720 363.670 399.005 ;
        RECT 364.510 395.720 365.510 399.005 ;
        RECT 366.350 395.720 367.350 399.005 ;
        RECT 368.190 395.720 368.730 399.005 ;
        RECT 369.570 395.720 370.570 399.005 ;
        RECT 371.410 395.720 372.410 399.005 ;
        RECT 373.250 395.720 374.250 399.005 ;
        RECT 375.090 395.720 376.090 399.005 ;
        RECT 376.930 395.720 377.470 399.005 ;
        RECT 378.310 395.720 379.310 399.005 ;
        RECT 380.150 395.720 381.150 399.005 ;
        RECT 381.990 395.720 382.990 399.005 ;
        RECT 383.830 395.720 384.370 399.005 ;
        RECT 385.210 395.720 386.210 399.005 ;
        RECT 387.050 395.720 388.050 399.005 ;
        RECT 388.890 395.720 389.890 399.005 ;
        RECT 390.730 395.720 391.730 399.005 ;
        RECT 392.570 395.720 393.110 399.005 ;
        RECT 393.950 395.720 394.950 399.005 ;
        RECT 395.790 395.720 396.790 399.005 ;
        RECT 397.630 395.720 398.630 399.005 ;
        RECT 0.560 4.280 399.180 395.720 ;
        RECT 1.110 0.835 1.650 4.280 ;
        RECT 2.490 0.835 3.490 4.280 ;
        RECT 4.330 0.835 4.870 4.280 ;
        RECT 5.710 0.835 6.710 4.280 ;
        RECT 7.550 0.835 8.550 4.280 ;
        RECT 9.390 0.835 9.930 4.280 ;
        RECT 10.770 0.835 11.770 4.280 ;
        RECT 12.610 0.835 13.610 4.280 ;
        RECT 14.450 0.835 14.990 4.280 ;
        RECT 15.830 0.835 16.830 4.280 ;
        RECT 17.670 0.835 18.670 4.280 ;
        RECT 19.510 0.835 20.050 4.280 ;
        RECT 20.890 0.835 21.890 4.280 ;
        RECT 22.730 0.835 23.730 4.280 ;
        RECT 24.570 0.835 25.110 4.280 ;
        RECT 25.950 0.835 26.950 4.280 ;
        RECT 27.790 0.835 28.790 4.280 ;
        RECT 29.630 0.835 30.170 4.280 ;
        RECT 31.010 0.835 32.010 4.280 ;
        RECT 32.850 0.835 33.850 4.280 ;
        RECT 34.690 0.835 35.230 4.280 ;
        RECT 36.070 0.835 37.070 4.280 ;
        RECT 37.910 0.835 38.910 4.280 ;
        RECT 39.750 0.835 40.290 4.280 ;
        RECT 41.130 0.835 42.130 4.280 ;
        RECT 42.970 0.835 43.970 4.280 ;
        RECT 44.810 0.835 45.350 4.280 ;
        RECT 46.190 0.835 47.190 4.280 ;
        RECT 48.030 0.835 49.030 4.280 ;
        RECT 49.870 0.835 50.410 4.280 ;
        RECT 51.250 0.835 52.250 4.280 ;
        RECT 53.090 0.835 53.630 4.280 ;
        RECT 54.470 0.835 55.470 4.280 ;
        RECT 56.310 0.835 57.310 4.280 ;
        RECT 58.150 0.835 58.690 4.280 ;
        RECT 59.530 0.835 60.530 4.280 ;
        RECT 61.370 0.835 62.370 4.280 ;
        RECT 63.210 0.835 63.750 4.280 ;
        RECT 64.590 0.835 65.590 4.280 ;
        RECT 66.430 0.835 67.430 4.280 ;
        RECT 68.270 0.835 68.810 4.280 ;
        RECT 69.650 0.835 70.650 4.280 ;
        RECT 71.490 0.835 72.490 4.280 ;
        RECT 73.330 0.835 73.870 4.280 ;
        RECT 74.710 0.835 75.710 4.280 ;
        RECT 76.550 0.835 77.550 4.280 ;
        RECT 78.390 0.835 78.930 4.280 ;
        RECT 79.770 0.835 80.770 4.280 ;
        RECT 81.610 0.835 82.610 4.280 ;
        RECT 83.450 0.835 83.990 4.280 ;
        RECT 84.830 0.835 85.830 4.280 ;
        RECT 86.670 0.835 87.670 4.280 ;
        RECT 88.510 0.835 89.050 4.280 ;
        RECT 89.890 0.835 90.890 4.280 ;
        RECT 91.730 0.835 92.730 4.280 ;
        RECT 93.570 0.835 94.110 4.280 ;
        RECT 94.950 0.835 95.950 4.280 ;
        RECT 96.790 0.835 97.790 4.280 ;
        RECT 98.630 0.835 99.170 4.280 ;
        RECT 100.010 0.835 101.010 4.280 ;
        RECT 101.850 0.835 102.390 4.280 ;
        RECT 103.230 0.835 104.230 4.280 ;
        RECT 105.070 0.835 106.070 4.280 ;
        RECT 106.910 0.835 107.450 4.280 ;
        RECT 108.290 0.835 109.290 4.280 ;
        RECT 110.130 0.835 111.130 4.280 ;
        RECT 111.970 0.835 112.510 4.280 ;
        RECT 113.350 0.835 114.350 4.280 ;
        RECT 115.190 0.835 116.190 4.280 ;
        RECT 117.030 0.835 117.570 4.280 ;
        RECT 118.410 0.835 119.410 4.280 ;
        RECT 120.250 0.835 121.250 4.280 ;
        RECT 122.090 0.835 122.630 4.280 ;
        RECT 123.470 0.835 124.470 4.280 ;
        RECT 125.310 0.835 126.310 4.280 ;
        RECT 127.150 0.835 127.690 4.280 ;
        RECT 128.530 0.835 129.530 4.280 ;
        RECT 130.370 0.835 131.370 4.280 ;
        RECT 132.210 0.835 132.750 4.280 ;
        RECT 133.590 0.835 134.590 4.280 ;
        RECT 135.430 0.835 136.430 4.280 ;
        RECT 137.270 0.835 137.810 4.280 ;
        RECT 138.650 0.835 139.650 4.280 ;
        RECT 140.490 0.835 141.490 4.280 ;
        RECT 142.330 0.835 142.870 4.280 ;
        RECT 143.710 0.835 144.710 4.280 ;
        RECT 145.550 0.835 146.550 4.280 ;
        RECT 147.390 0.835 147.930 4.280 ;
        RECT 148.770 0.835 149.770 4.280 ;
        RECT 150.610 0.835 151.150 4.280 ;
        RECT 151.990 0.835 152.990 4.280 ;
        RECT 153.830 0.835 154.830 4.280 ;
        RECT 155.670 0.835 156.210 4.280 ;
        RECT 157.050 0.835 158.050 4.280 ;
        RECT 158.890 0.835 159.890 4.280 ;
        RECT 160.730 0.835 161.270 4.280 ;
        RECT 162.110 0.835 163.110 4.280 ;
        RECT 163.950 0.835 164.950 4.280 ;
        RECT 165.790 0.835 166.330 4.280 ;
        RECT 167.170 0.835 168.170 4.280 ;
        RECT 169.010 0.835 170.010 4.280 ;
        RECT 170.850 0.835 171.390 4.280 ;
        RECT 172.230 0.835 173.230 4.280 ;
        RECT 174.070 0.835 175.070 4.280 ;
        RECT 175.910 0.835 176.450 4.280 ;
        RECT 177.290 0.835 178.290 4.280 ;
        RECT 179.130 0.835 180.130 4.280 ;
        RECT 180.970 0.835 181.510 4.280 ;
        RECT 182.350 0.835 183.350 4.280 ;
        RECT 184.190 0.835 185.190 4.280 ;
        RECT 186.030 0.835 186.570 4.280 ;
        RECT 187.410 0.835 188.410 4.280 ;
        RECT 189.250 0.835 190.250 4.280 ;
        RECT 191.090 0.835 191.630 4.280 ;
        RECT 192.470 0.835 193.470 4.280 ;
        RECT 194.310 0.835 195.310 4.280 ;
        RECT 196.150 0.835 196.690 4.280 ;
        RECT 197.530 0.835 198.530 4.280 ;
        RECT 199.370 0.835 200.370 4.280 ;
        RECT 201.210 0.835 201.750 4.280 ;
        RECT 202.590 0.835 203.590 4.280 ;
        RECT 204.430 0.835 204.970 4.280 ;
        RECT 205.810 0.835 206.810 4.280 ;
        RECT 207.650 0.835 208.650 4.280 ;
        RECT 209.490 0.835 210.030 4.280 ;
        RECT 210.870 0.835 211.870 4.280 ;
        RECT 212.710 0.835 213.710 4.280 ;
        RECT 214.550 0.835 215.090 4.280 ;
        RECT 215.930 0.835 216.930 4.280 ;
        RECT 217.770 0.835 218.770 4.280 ;
        RECT 219.610 0.835 220.150 4.280 ;
        RECT 220.990 0.835 221.990 4.280 ;
        RECT 222.830 0.835 223.830 4.280 ;
        RECT 224.670 0.835 225.210 4.280 ;
        RECT 226.050 0.835 227.050 4.280 ;
        RECT 227.890 0.835 228.890 4.280 ;
        RECT 229.730 0.835 230.270 4.280 ;
        RECT 231.110 0.835 232.110 4.280 ;
        RECT 232.950 0.835 233.950 4.280 ;
        RECT 234.790 0.835 235.330 4.280 ;
        RECT 236.170 0.835 237.170 4.280 ;
        RECT 238.010 0.835 239.010 4.280 ;
        RECT 239.850 0.835 240.390 4.280 ;
        RECT 241.230 0.835 242.230 4.280 ;
        RECT 243.070 0.835 244.070 4.280 ;
        RECT 244.910 0.835 245.450 4.280 ;
        RECT 246.290 0.835 247.290 4.280 ;
        RECT 248.130 0.835 249.130 4.280 ;
        RECT 249.970 0.835 250.510 4.280 ;
        RECT 251.350 0.835 252.350 4.280 ;
        RECT 253.190 0.835 253.730 4.280 ;
        RECT 254.570 0.835 255.570 4.280 ;
        RECT 256.410 0.835 257.410 4.280 ;
        RECT 258.250 0.835 258.790 4.280 ;
        RECT 259.630 0.835 260.630 4.280 ;
        RECT 261.470 0.835 262.470 4.280 ;
        RECT 263.310 0.835 263.850 4.280 ;
        RECT 264.690 0.835 265.690 4.280 ;
        RECT 266.530 0.835 267.530 4.280 ;
        RECT 268.370 0.835 268.910 4.280 ;
        RECT 269.750 0.835 270.750 4.280 ;
        RECT 271.590 0.835 272.590 4.280 ;
        RECT 273.430 0.835 273.970 4.280 ;
        RECT 274.810 0.835 275.810 4.280 ;
        RECT 276.650 0.835 277.650 4.280 ;
        RECT 278.490 0.835 279.030 4.280 ;
        RECT 279.870 0.835 280.870 4.280 ;
        RECT 281.710 0.835 282.710 4.280 ;
        RECT 283.550 0.835 284.090 4.280 ;
        RECT 284.930 0.835 285.930 4.280 ;
        RECT 286.770 0.835 287.770 4.280 ;
        RECT 288.610 0.835 289.150 4.280 ;
        RECT 289.990 0.835 290.990 4.280 ;
        RECT 291.830 0.835 292.830 4.280 ;
        RECT 293.670 0.835 294.210 4.280 ;
        RECT 295.050 0.835 296.050 4.280 ;
        RECT 296.890 0.835 297.890 4.280 ;
        RECT 298.730 0.835 299.270 4.280 ;
        RECT 300.110 0.835 301.110 4.280 ;
        RECT 301.950 0.835 302.490 4.280 ;
        RECT 303.330 0.835 304.330 4.280 ;
        RECT 305.170 0.835 306.170 4.280 ;
        RECT 307.010 0.835 307.550 4.280 ;
        RECT 308.390 0.835 309.390 4.280 ;
        RECT 310.230 0.835 311.230 4.280 ;
        RECT 312.070 0.835 312.610 4.280 ;
        RECT 313.450 0.835 314.450 4.280 ;
        RECT 315.290 0.835 316.290 4.280 ;
        RECT 317.130 0.835 317.670 4.280 ;
        RECT 318.510 0.835 319.510 4.280 ;
        RECT 320.350 0.835 321.350 4.280 ;
        RECT 322.190 0.835 322.730 4.280 ;
        RECT 323.570 0.835 324.570 4.280 ;
        RECT 325.410 0.835 326.410 4.280 ;
        RECT 327.250 0.835 327.790 4.280 ;
        RECT 328.630 0.835 329.630 4.280 ;
        RECT 330.470 0.835 331.470 4.280 ;
        RECT 332.310 0.835 332.850 4.280 ;
        RECT 333.690 0.835 334.690 4.280 ;
        RECT 335.530 0.835 336.530 4.280 ;
        RECT 337.370 0.835 337.910 4.280 ;
        RECT 338.750 0.835 339.750 4.280 ;
        RECT 340.590 0.835 341.590 4.280 ;
        RECT 342.430 0.835 342.970 4.280 ;
        RECT 343.810 0.835 344.810 4.280 ;
        RECT 345.650 0.835 346.650 4.280 ;
        RECT 347.490 0.835 348.030 4.280 ;
        RECT 348.870 0.835 349.870 4.280 ;
        RECT 350.710 0.835 351.250 4.280 ;
        RECT 352.090 0.835 353.090 4.280 ;
        RECT 353.930 0.835 354.930 4.280 ;
        RECT 355.770 0.835 356.310 4.280 ;
        RECT 357.150 0.835 358.150 4.280 ;
        RECT 358.990 0.835 359.990 4.280 ;
        RECT 360.830 0.835 361.370 4.280 ;
        RECT 362.210 0.835 363.210 4.280 ;
        RECT 364.050 0.835 365.050 4.280 ;
        RECT 365.890 0.835 366.430 4.280 ;
        RECT 367.270 0.835 368.270 4.280 ;
        RECT 369.110 0.835 370.110 4.280 ;
        RECT 370.950 0.835 371.490 4.280 ;
        RECT 372.330 0.835 373.330 4.280 ;
        RECT 374.170 0.835 375.170 4.280 ;
        RECT 376.010 0.835 376.550 4.280 ;
        RECT 377.390 0.835 378.390 4.280 ;
        RECT 379.230 0.835 380.230 4.280 ;
        RECT 381.070 0.835 381.610 4.280 ;
        RECT 382.450 0.835 383.450 4.280 ;
        RECT 384.290 0.835 385.290 4.280 ;
        RECT 386.130 0.835 386.670 4.280 ;
        RECT 387.510 0.835 388.510 4.280 ;
        RECT 389.350 0.835 390.350 4.280 ;
        RECT 391.190 0.835 391.730 4.280 ;
        RECT 392.570 0.835 393.570 4.280 ;
        RECT 394.410 0.835 395.410 4.280 ;
        RECT 396.250 0.835 396.790 4.280 ;
        RECT 397.630 0.835 398.630 4.280 ;
      LAYER met3 ;
        RECT 4.400 398.120 395.600 398.985 ;
        RECT 4.000 397.480 395.600 398.120 ;
        RECT 4.400 396.080 395.600 397.480 ;
        RECT 4.000 395.440 395.600 396.080 ;
        RECT 4.400 395.400 395.600 395.440 ;
        RECT 4.400 394.760 396.000 395.400 ;
        RECT 4.400 392.680 395.600 394.760 ;
        RECT 4.000 392.040 395.600 392.680 ;
        RECT 4.400 390.640 395.600 392.040 ;
        RECT 4.000 390.000 396.000 390.640 ;
        RECT 4.400 387.240 395.600 390.000 ;
        RECT 4.000 386.600 395.600 387.240 ;
        RECT 4.400 385.880 395.600 386.600 ;
        RECT 4.400 385.240 396.000 385.880 ;
        RECT 4.400 385.200 395.600 385.240 ;
        RECT 4.000 384.560 395.600 385.200 ;
        RECT 4.400 381.800 395.600 384.560 ;
        RECT 4.000 381.160 395.600 381.800 ;
        RECT 4.400 381.120 395.600 381.160 ;
        RECT 4.400 380.480 396.000 381.120 ;
        RECT 4.400 379.760 395.600 380.480 ;
        RECT 4.000 379.120 395.600 379.760 ;
        RECT 4.400 376.360 395.600 379.120 ;
        RECT 4.000 375.720 396.000 376.360 ;
        RECT 4.400 374.320 395.600 375.720 ;
        RECT 4.000 373.680 395.600 374.320 ;
        RECT 4.400 370.920 395.600 373.680 ;
        RECT 4.000 370.280 395.600 370.920 ;
        RECT 4.400 370.240 395.600 370.280 ;
        RECT 4.400 369.600 396.000 370.240 ;
        RECT 4.400 368.880 395.600 369.600 ;
        RECT 4.000 368.240 395.600 368.880 ;
        RECT 4.400 365.480 395.600 368.240 ;
        RECT 4.000 364.840 396.000 365.480 ;
        RECT 4.400 363.440 395.600 364.840 ;
        RECT 4.000 362.800 395.600 363.440 ;
        RECT 4.400 360.720 395.600 362.800 ;
        RECT 4.400 360.080 396.000 360.720 ;
        RECT 4.400 360.040 395.600 360.080 ;
        RECT 4.000 359.400 395.600 360.040 ;
        RECT 4.400 358.000 395.600 359.400 ;
        RECT 4.000 357.360 395.600 358.000 ;
        RECT 4.400 355.960 395.600 357.360 ;
        RECT 4.400 355.320 396.000 355.960 ;
        RECT 4.400 354.600 395.600 355.320 ;
        RECT 4.000 353.960 395.600 354.600 ;
        RECT 4.400 352.560 395.600 353.960 ;
        RECT 4.000 351.920 395.600 352.560 ;
        RECT 4.400 351.200 395.600 351.920 ;
        RECT 4.400 350.560 396.000 351.200 ;
        RECT 4.400 349.160 395.600 350.560 ;
        RECT 4.000 348.520 395.600 349.160 ;
        RECT 4.400 347.120 395.600 348.520 ;
        RECT 4.000 346.480 395.600 347.120 ;
        RECT 4.400 346.440 395.600 346.480 ;
        RECT 4.400 345.800 396.000 346.440 ;
        RECT 4.400 343.720 395.600 345.800 ;
        RECT 4.000 343.080 395.600 343.720 ;
        RECT 4.400 341.680 395.600 343.080 ;
        RECT 4.000 341.040 395.600 341.680 ;
        RECT 4.400 340.320 395.600 341.040 ;
        RECT 4.400 339.680 396.000 340.320 ;
        RECT 4.400 338.280 395.600 339.680 ;
        RECT 4.000 337.640 395.600 338.280 ;
        RECT 4.400 336.240 395.600 337.640 ;
        RECT 4.000 335.600 395.600 336.240 ;
        RECT 4.400 335.560 395.600 335.600 ;
        RECT 4.400 334.920 396.000 335.560 ;
        RECT 4.400 332.840 395.600 334.920 ;
        RECT 4.000 332.200 395.600 332.840 ;
        RECT 4.400 330.800 395.600 332.200 ;
        RECT 4.000 330.160 396.000 330.800 ;
        RECT 4.400 327.400 395.600 330.160 ;
        RECT 4.000 326.760 395.600 327.400 ;
        RECT 4.400 326.040 395.600 326.760 ;
        RECT 4.400 325.400 396.000 326.040 ;
        RECT 4.400 325.360 395.600 325.400 ;
        RECT 4.000 324.720 395.600 325.360 ;
        RECT 4.400 321.960 395.600 324.720 ;
        RECT 4.000 321.320 395.600 321.960 ;
        RECT 4.400 321.280 395.600 321.320 ;
        RECT 4.400 320.640 396.000 321.280 ;
        RECT 4.400 319.920 395.600 320.640 ;
        RECT 4.000 319.280 395.600 319.920 ;
        RECT 4.400 316.520 395.600 319.280 ;
        RECT 4.000 315.880 396.000 316.520 ;
        RECT 4.400 314.480 395.600 315.880 ;
        RECT 4.000 313.840 395.600 314.480 ;
        RECT 4.400 311.080 395.600 313.840 ;
        RECT 4.000 310.440 395.600 311.080 ;
        RECT 4.400 310.400 395.600 310.440 ;
        RECT 4.400 309.760 396.000 310.400 ;
        RECT 4.400 309.040 395.600 309.760 ;
        RECT 4.000 308.400 395.600 309.040 ;
        RECT 4.400 305.640 395.600 308.400 ;
        RECT 4.000 305.000 396.000 305.640 ;
        RECT 4.400 303.600 395.600 305.000 ;
        RECT 4.000 302.960 395.600 303.600 ;
        RECT 4.400 300.880 395.600 302.960 ;
        RECT 4.400 300.240 396.000 300.880 ;
        RECT 4.400 300.200 395.600 300.240 ;
        RECT 4.000 299.560 395.600 300.200 ;
        RECT 4.400 298.160 395.600 299.560 ;
        RECT 4.000 297.520 395.600 298.160 ;
        RECT 4.400 296.120 395.600 297.520 ;
        RECT 4.000 295.480 396.000 296.120 ;
        RECT 4.400 292.720 395.600 295.480 ;
        RECT 4.000 292.080 395.600 292.720 ;
        RECT 4.400 291.360 395.600 292.080 ;
        RECT 4.400 290.720 396.000 291.360 ;
        RECT 4.400 290.680 395.600 290.720 ;
        RECT 4.000 290.040 395.600 290.680 ;
        RECT 4.400 287.280 395.600 290.040 ;
        RECT 4.000 286.640 395.600 287.280 ;
        RECT 4.400 285.240 395.600 286.640 ;
        RECT 4.000 284.600 396.000 285.240 ;
        RECT 4.400 281.840 395.600 284.600 ;
        RECT 4.000 281.200 395.600 281.840 ;
        RECT 4.400 280.480 395.600 281.200 ;
        RECT 4.400 279.840 396.000 280.480 ;
        RECT 4.400 279.800 395.600 279.840 ;
        RECT 4.000 279.160 395.600 279.800 ;
        RECT 4.400 276.400 395.600 279.160 ;
        RECT 4.000 275.760 395.600 276.400 ;
        RECT 4.400 275.720 395.600 275.760 ;
        RECT 4.400 275.080 396.000 275.720 ;
        RECT 4.400 274.360 395.600 275.080 ;
        RECT 4.000 273.720 395.600 274.360 ;
        RECT 4.400 270.960 395.600 273.720 ;
        RECT 4.000 270.320 396.000 270.960 ;
        RECT 4.400 268.920 395.600 270.320 ;
        RECT 4.000 268.280 395.600 268.920 ;
        RECT 4.400 266.200 395.600 268.280 ;
        RECT 4.400 265.560 396.000 266.200 ;
        RECT 4.400 265.520 395.600 265.560 ;
        RECT 4.000 264.880 395.600 265.520 ;
        RECT 4.400 263.480 395.600 264.880 ;
        RECT 4.000 262.840 395.600 263.480 ;
        RECT 4.400 261.440 395.600 262.840 ;
        RECT 4.400 260.800 396.000 261.440 ;
        RECT 4.400 260.080 395.600 260.800 ;
        RECT 4.000 259.440 395.600 260.080 ;
        RECT 4.400 258.040 395.600 259.440 ;
        RECT 4.000 257.400 395.600 258.040 ;
        RECT 4.400 255.320 395.600 257.400 ;
        RECT 4.400 254.680 396.000 255.320 ;
        RECT 4.400 254.640 395.600 254.680 ;
        RECT 4.000 254.000 395.600 254.640 ;
        RECT 4.400 252.600 395.600 254.000 ;
        RECT 4.000 251.960 395.600 252.600 ;
        RECT 4.400 250.560 395.600 251.960 ;
        RECT 4.400 249.920 396.000 250.560 ;
        RECT 4.400 249.200 395.600 249.920 ;
        RECT 4.000 248.560 395.600 249.200 ;
        RECT 4.400 247.160 395.600 248.560 ;
        RECT 4.000 246.520 395.600 247.160 ;
        RECT 4.400 245.800 395.600 246.520 ;
        RECT 4.400 245.160 396.000 245.800 ;
        RECT 4.400 243.760 395.600 245.160 ;
        RECT 4.000 243.120 395.600 243.760 ;
        RECT 4.400 241.720 395.600 243.120 ;
        RECT 4.000 241.080 395.600 241.720 ;
        RECT 4.400 241.040 395.600 241.080 ;
        RECT 4.400 240.400 396.000 241.040 ;
        RECT 4.400 238.320 395.600 240.400 ;
        RECT 4.000 237.680 395.600 238.320 ;
        RECT 4.400 236.280 395.600 237.680 ;
        RECT 4.000 235.640 396.000 236.280 ;
        RECT 4.400 232.880 395.600 235.640 ;
        RECT 4.000 232.240 395.600 232.880 ;
        RECT 4.400 231.520 395.600 232.240 ;
        RECT 4.400 230.880 396.000 231.520 ;
        RECT 4.400 230.840 395.600 230.880 ;
        RECT 4.000 230.200 395.600 230.840 ;
        RECT 4.400 227.440 395.600 230.200 ;
        RECT 4.000 226.800 395.600 227.440 ;
        RECT 4.400 225.400 395.600 226.800 ;
        RECT 4.000 224.760 396.000 225.400 ;
        RECT 4.400 222.000 395.600 224.760 ;
        RECT 4.000 221.360 395.600 222.000 ;
        RECT 4.400 220.640 395.600 221.360 ;
        RECT 4.400 220.000 396.000 220.640 ;
        RECT 4.400 219.960 395.600 220.000 ;
        RECT 4.000 219.320 395.600 219.960 ;
        RECT 4.400 216.560 395.600 219.320 ;
        RECT 4.000 215.920 395.600 216.560 ;
        RECT 4.400 215.880 395.600 215.920 ;
        RECT 4.400 215.240 396.000 215.880 ;
        RECT 4.400 214.520 395.600 215.240 ;
        RECT 4.000 213.880 395.600 214.520 ;
        RECT 4.400 211.120 395.600 213.880 ;
        RECT 4.000 210.480 396.000 211.120 ;
        RECT 4.400 209.080 395.600 210.480 ;
        RECT 4.000 208.440 395.600 209.080 ;
        RECT 4.400 206.360 395.600 208.440 ;
        RECT 4.400 205.720 396.000 206.360 ;
        RECT 4.400 205.680 395.600 205.720 ;
        RECT 4.000 205.040 395.600 205.680 ;
        RECT 4.400 203.640 395.600 205.040 ;
        RECT 4.000 203.000 395.600 203.640 ;
        RECT 4.400 200.240 395.600 203.000 ;
        RECT 4.000 199.600 396.000 200.240 ;
        RECT 4.400 198.200 395.600 199.600 ;
        RECT 4.000 197.560 395.600 198.200 ;
        RECT 4.400 196.160 395.600 197.560 ;
        RECT 4.000 195.520 395.600 196.160 ;
        RECT 4.400 195.480 395.600 195.520 ;
        RECT 4.400 194.840 396.000 195.480 ;
        RECT 4.400 192.760 395.600 194.840 ;
        RECT 4.000 192.120 395.600 192.760 ;
        RECT 4.400 190.720 395.600 192.120 ;
        RECT 4.000 190.080 396.000 190.720 ;
        RECT 4.400 187.320 395.600 190.080 ;
        RECT 4.000 186.680 395.600 187.320 ;
        RECT 4.400 185.960 395.600 186.680 ;
        RECT 4.400 185.320 396.000 185.960 ;
        RECT 4.400 185.280 395.600 185.320 ;
        RECT 4.000 184.640 395.600 185.280 ;
        RECT 4.400 181.880 395.600 184.640 ;
        RECT 4.000 181.240 395.600 181.880 ;
        RECT 4.400 181.200 395.600 181.240 ;
        RECT 4.400 180.560 396.000 181.200 ;
        RECT 4.400 179.840 395.600 180.560 ;
        RECT 4.000 179.200 395.600 179.840 ;
        RECT 4.400 176.440 395.600 179.200 ;
        RECT 4.000 175.800 396.000 176.440 ;
        RECT 4.400 174.400 395.600 175.800 ;
        RECT 4.000 173.760 395.600 174.400 ;
        RECT 4.400 171.000 395.600 173.760 ;
        RECT 4.000 170.360 395.600 171.000 ;
        RECT 4.400 170.320 395.600 170.360 ;
        RECT 4.400 169.680 396.000 170.320 ;
        RECT 4.400 168.960 395.600 169.680 ;
        RECT 4.000 168.320 395.600 168.960 ;
        RECT 4.400 165.560 395.600 168.320 ;
        RECT 4.000 164.920 396.000 165.560 ;
        RECT 4.400 163.520 395.600 164.920 ;
        RECT 4.000 162.880 395.600 163.520 ;
        RECT 4.400 160.800 395.600 162.880 ;
        RECT 4.400 160.160 396.000 160.800 ;
        RECT 4.400 160.120 395.600 160.160 ;
        RECT 4.000 159.480 395.600 160.120 ;
        RECT 4.400 158.080 395.600 159.480 ;
        RECT 4.000 157.440 395.600 158.080 ;
        RECT 4.400 156.040 395.600 157.440 ;
        RECT 4.400 155.400 396.000 156.040 ;
        RECT 4.400 154.680 395.600 155.400 ;
        RECT 4.000 154.040 395.600 154.680 ;
        RECT 4.400 152.640 395.600 154.040 ;
        RECT 4.000 152.000 395.600 152.640 ;
        RECT 4.400 151.280 395.600 152.000 ;
        RECT 4.400 150.640 396.000 151.280 ;
        RECT 4.400 149.240 395.600 150.640 ;
        RECT 4.000 148.600 395.600 149.240 ;
        RECT 4.400 147.200 395.600 148.600 ;
        RECT 4.000 146.560 395.600 147.200 ;
        RECT 4.400 146.520 395.600 146.560 ;
        RECT 4.400 145.880 396.000 146.520 ;
        RECT 4.400 143.800 395.600 145.880 ;
        RECT 4.000 143.160 395.600 143.800 ;
        RECT 4.400 141.760 395.600 143.160 ;
        RECT 4.000 141.120 395.600 141.760 ;
        RECT 4.400 140.400 395.600 141.120 ;
        RECT 4.400 139.760 396.000 140.400 ;
        RECT 4.400 138.360 395.600 139.760 ;
        RECT 4.000 137.720 395.600 138.360 ;
        RECT 4.400 136.320 395.600 137.720 ;
        RECT 4.000 135.680 395.600 136.320 ;
        RECT 4.400 135.640 395.600 135.680 ;
        RECT 4.400 135.000 396.000 135.640 ;
        RECT 4.400 132.920 395.600 135.000 ;
        RECT 4.000 132.280 395.600 132.920 ;
        RECT 4.400 130.880 395.600 132.280 ;
        RECT 4.000 130.240 396.000 130.880 ;
        RECT 4.400 127.480 395.600 130.240 ;
        RECT 4.000 126.840 395.600 127.480 ;
        RECT 4.400 126.120 395.600 126.840 ;
        RECT 4.400 125.480 396.000 126.120 ;
        RECT 4.400 125.440 395.600 125.480 ;
        RECT 4.000 124.800 395.600 125.440 ;
        RECT 4.400 122.040 395.600 124.800 ;
        RECT 4.000 121.400 395.600 122.040 ;
        RECT 4.400 121.360 395.600 121.400 ;
        RECT 4.400 120.720 396.000 121.360 ;
        RECT 4.400 120.000 395.600 120.720 ;
        RECT 4.000 119.360 395.600 120.000 ;
        RECT 4.400 116.600 395.600 119.360 ;
        RECT 4.000 115.960 396.000 116.600 ;
        RECT 4.400 114.560 395.600 115.960 ;
        RECT 4.000 113.920 395.600 114.560 ;
        RECT 4.400 111.160 395.600 113.920 ;
        RECT 4.000 110.520 395.600 111.160 ;
        RECT 4.400 110.480 395.600 110.520 ;
        RECT 4.400 109.840 396.000 110.480 ;
        RECT 4.400 109.120 395.600 109.840 ;
        RECT 4.000 108.480 395.600 109.120 ;
        RECT 4.400 105.720 395.600 108.480 ;
        RECT 4.000 105.080 396.000 105.720 ;
        RECT 4.400 103.680 395.600 105.080 ;
        RECT 4.000 103.040 395.600 103.680 ;
        RECT 4.400 100.960 395.600 103.040 ;
        RECT 4.400 100.320 396.000 100.960 ;
        RECT 4.400 100.280 395.600 100.320 ;
        RECT 4.000 99.640 395.600 100.280 ;
        RECT 4.400 98.240 395.600 99.640 ;
        RECT 4.000 97.600 395.600 98.240 ;
        RECT 4.400 96.200 395.600 97.600 ;
        RECT 4.000 95.560 396.000 96.200 ;
        RECT 4.400 92.800 395.600 95.560 ;
        RECT 4.000 92.160 395.600 92.800 ;
        RECT 4.400 91.440 395.600 92.160 ;
        RECT 4.400 90.800 396.000 91.440 ;
        RECT 4.400 90.760 395.600 90.800 ;
        RECT 4.000 90.120 395.600 90.760 ;
        RECT 4.400 87.360 395.600 90.120 ;
        RECT 4.000 86.720 395.600 87.360 ;
        RECT 4.400 85.320 395.600 86.720 ;
        RECT 4.000 84.680 396.000 85.320 ;
        RECT 4.400 81.920 395.600 84.680 ;
        RECT 4.000 81.280 395.600 81.920 ;
        RECT 4.400 80.560 395.600 81.280 ;
        RECT 4.400 79.920 396.000 80.560 ;
        RECT 4.400 79.880 395.600 79.920 ;
        RECT 4.000 79.240 395.600 79.880 ;
        RECT 4.400 76.480 395.600 79.240 ;
        RECT 4.000 75.840 395.600 76.480 ;
        RECT 4.400 75.800 395.600 75.840 ;
        RECT 4.400 75.160 396.000 75.800 ;
        RECT 4.400 74.440 395.600 75.160 ;
        RECT 4.000 73.800 395.600 74.440 ;
        RECT 4.400 71.040 395.600 73.800 ;
        RECT 4.000 70.400 396.000 71.040 ;
        RECT 4.400 69.000 395.600 70.400 ;
        RECT 4.000 68.360 395.600 69.000 ;
        RECT 4.400 66.280 395.600 68.360 ;
        RECT 4.400 65.640 396.000 66.280 ;
        RECT 4.400 65.600 395.600 65.640 ;
        RECT 4.000 64.960 395.600 65.600 ;
        RECT 4.400 63.560 395.600 64.960 ;
        RECT 4.000 62.920 395.600 63.560 ;
        RECT 4.400 61.520 395.600 62.920 ;
        RECT 4.400 60.880 396.000 61.520 ;
        RECT 4.400 60.160 395.600 60.880 ;
        RECT 4.000 59.520 395.600 60.160 ;
        RECT 4.400 58.120 395.600 59.520 ;
        RECT 4.000 57.480 395.600 58.120 ;
        RECT 4.400 55.400 395.600 57.480 ;
        RECT 4.400 54.760 396.000 55.400 ;
        RECT 4.400 54.720 395.600 54.760 ;
        RECT 4.000 54.080 395.600 54.720 ;
        RECT 4.400 52.680 395.600 54.080 ;
        RECT 4.000 52.040 395.600 52.680 ;
        RECT 4.400 50.640 395.600 52.040 ;
        RECT 4.400 50.000 396.000 50.640 ;
        RECT 4.400 49.280 395.600 50.000 ;
        RECT 4.000 48.640 395.600 49.280 ;
        RECT 4.400 47.240 395.600 48.640 ;
        RECT 4.000 46.600 395.600 47.240 ;
        RECT 4.400 45.880 395.600 46.600 ;
        RECT 4.400 45.240 396.000 45.880 ;
        RECT 4.400 43.840 395.600 45.240 ;
        RECT 4.000 43.200 395.600 43.840 ;
        RECT 4.400 41.800 395.600 43.200 ;
        RECT 4.000 41.160 395.600 41.800 ;
        RECT 4.400 41.120 395.600 41.160 ;
        RECT 4.400 40.480 396.000 41.120 ;
        RECT 4.400 38.400 395.600 40.480 ;
        RECT 4.000 37.760 395.600 38.400 ;
        RECT 4.400 36.360 395.600 37.760 ;
        RECT 4.000 35.720 396.000 36.360 ;
        RECT 4.400 32.960 395.600 35.720 ;
        RECT 4.000 32.320 395.600 32.960 ;
        RECT 4.400 31.600 395.600 32.320 ;
        RECT 4.400 30.960 396.000 31.600 ;
        RECT 4.400 30.920 395.600 30.960 ;
        RECT 4.000 30.280 395.600 30.920 ;
        RECT 4.400 27.520 395.600 30.280 ;
        RECT 4.000 26.880 395.600 27.520 ;
        RECT 4.400 25.480 395.600 26.880 ;
        RECT 4.000 24.840 396.000 25.480 ;
        RECT 4.400 22.080 395.600 24.840 ;
        RECT 4.000 21.440 395.600 22.080 ;
        RECT 4.400 20.720 395.600 21.440 ;
        RECT 4.400 20.080 396.000 20.720 ;
        RECT 4.400 20.040 395.600 20.080 ;
        RECT 4.000 19.400 395.600 20.040 ;
        RECT 4.400 16.640 395.600 19.400 ;
        RECT 4.000 16.000 395.600 16.640 ;
        RECT 4.400 15.960 395.600 16.000 ;
        RECT 4.400 15.320 396.000 15.960 ;
        RECT 4.400 14.600 395.600 15.320 ;
        RECT 4.000 13.960 395.600 14.600 ;
        RECT 4.400 11.200 395.600 13.960 ;
        RECT 4.000 10.560 396.000 11.200 ;
        RECT 4.400 9.160 395.600 10.560 ;
        RECT 4.000 8.520 395.600 9.160 ;
        RECT 4.400 6.440 395.600 8.520 ;
        RECT 4.400 5.800 396.000 6.440 ;
        RECT 4.400 5.760 395.600 5.800 ;
        RECT 4.000 5.120 395.600 5.760 ;
        RECT 4.400 3.720 395.600 5.120 ;
        RECT 4.000 3.080 395.600 3.720 ;
        RECT 4.400 0.855 395.600 3.080 ;
      LAYER met4 ;
        RECT 15.935 10.240 20.640 227.625 ;
        RECT 23.040 10.240 97.440 227.625 ;
        RECT 99.840 10.240 174.240 227.625 ;
        RECT 176.640 10.240 251.040 227.625 ;
        RECT 253.440 10.240 327.840 227.625 ;
        RECT 330.240 10.240 374.145 227.625 ;
        RECT 15.935 9.015 374.145 10.240 ;
  END
END chip_controller
END LIBRARY

