VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 23.160 1500.000 23.760 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.930 0.000 1244.210 4.000 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1311.760 1500.000 1312.360 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.350 0.000 1279.630 4.000 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1274.360 4.000 1274.960 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 1496.000 1274.110 1500.000 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1344.400 1500.000 1345.000 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 0.000 1314.590 4.000 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.770 1496.000 1292.050 1500.000 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 0.000 1350.010 4.000 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1307.680 4.000 1308.280 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1324.680 4.000 1325.280 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1341.000 4.000 1341.600 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1393.360 1500.000 1393.960 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 1496.000 1364.270 1500.000 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1409.680 1500.000 1410.280 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.270 1496.000 1418.550 1500.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.570 0.000 1420.850 4.000 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1358.000 4.000 1358.600 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.050 0.000 1438.330 4.000 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 1496.000 315.930 1500.000 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1442.320 1500.000 1442.920 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1458.640 1500.000 1459.240 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1491.280 1500.000 1491.880 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1424.640 4.000 1425.240 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 0.000 1491.230 4.000 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1457.960 4.000 1458.560 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1474.280 4.000 1474.880 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 1496.000 334.330 1500.000 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 333.240 1500.000 333.840 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 398.520 1500.000 399.120 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 1496.000 406.550 1500.000 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 1496.000 99.270 1500.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 480.120 1500.000 480.720 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 1496.000 496.710 1500.000 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 545.400 1500.000 546.000 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1496.000 550.990 1500.000 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 594.360 1500.000 594.960 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 643.320 1500.000 643.920 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 72.120 1500.000 72.720 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 0.000 732.230 4.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 724.920 1500.000 725.520 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 741.240 1500.000 741.840 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 1496.000 677.490 1500.000 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.920 4.000 708.520 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 757.560 1500.000 758.160 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 1496.000 695.430 1500.000 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 789.520 1500.000 790.120 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 1496.000 713.830 1500.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 0.000 873.450 4.000 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 1496.000 731.770 1500.000 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 0.000 891.390 4.000 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 1496.000 749.710 1500.000 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 1496.000 786.050 1500.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 774.560 4.000 775.160 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 1496.000 803.990 1500.000 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 887.440 1500.000 888.040 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 1496.000 822.390 1500.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.880 4.000 825.480 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 0.000 908.870 4.000 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 0.000 926.350 4.000 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 920.080 1500.000 920.680 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.430 0.000 979.710 4.000 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 137.400 1500.000 138.000 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 1496.000 876.210 1500.000 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 1496.000 894.610 1500.000 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 1496.000 912.550 1500.000 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 936.400 1500.000 937.000 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 1496.000 948.890 1500.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.160 4.000 958.760 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 952.720 1500.000 953.320 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 1496.000 984.770 1500.000 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 969.040 1500.000 969.640 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 170.040 1500.000 170.640 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.800 4.000 1025.400 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 985.360 1500.000 985.960 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1001.680 1500.000 1002.280 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 0.000 1085.510 4.000 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.130 0.000 1138.410 4.000 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.770 1496.000 1039.050 1500.000 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 1496.000 1075.390 1500.000 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1050.640 1500.000 1051.240 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1083.280 1500.000 1083.880 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 1496.000 1093.330 1500.000 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 1496.000 1111.270 1500.000 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.550 0.000 1173.830 4.000 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930 1496.000 1129.210 1500.000 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1115.920 1500.000 1116.520 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1158.080 4.000 1158.680 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 1496.000 1147.610 1500.000 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.270 1496.000 1165.550 1500.000 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1181.200 1500.000 1181.800 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1213.840 1500.000 1214.440 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.030 0.000 1191.310 4.000 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 0.000 1208.790 4.000 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1279.120 1500.000 1279.720 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1295.440 1500.000 1296.040 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 1496.000 1183.490 1500.000 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.720 4.000 1225.320 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.040 4.000 1241.640 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 1496.000 1219.830 1500.000 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 316.920 1500.000 317.520 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 349.560 1500.000 350.160 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 447.480 1500.000 448.080 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 463.800 1500.000 464.400 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1496.000 460.830 1500.000 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 1496.000 515.110 1500.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 561.720 1500.000 562.320 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 1496.000 587.330 1500.000 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 1496.000 207.830 1500.000 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 202.680 1500.000 203.280 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 1496.000 44.990 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 1496.000 81.330 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 7.520 1500.000 8.120 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 1496.000 62.930 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 251.640 1500.000 252.240 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 267.960 1500.000 268.560 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 1496.000 370.210 1500.000 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 382.200 1500.000 382.800 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 1496.000 388.610 1500.000 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 55.800 1500.000 56.400 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 88.440 1500.000 89.040 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 104.760 1500.000 105.360 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 1496.000 171.490 1500.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 186.360 1500.000 186.960 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 1496.000 225.770 1500.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 219.000 1500.000 219.600 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.490 1496.000 1237.770 1500.000 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.410 0.000 1261.690 4.000 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.430 1496.000 1255.710 1500.000 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1291.360 4.000 1291.960 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1328.080 1500.000 1328.680 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.830 0.000 1297.110 4.000 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.250 0.000 1332.530 4.000 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 1496.000 1309.990 1500.000 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.670 0.000 1367.950 4.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1360.720 1500.000 1361.320 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 1496.000 280.050 1500.000 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.110 1496.000 1328.390 1500.000 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1377.040 1500.000 1377.640 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 1496.000 1346.330 1500.000 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.630 0.000 1402.910 4.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 1496.000 1382.210 1500.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.330 1496.000 1400.610 1500.000 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 1496.000 1436.490 1500.000 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1426.000 1500.000 1426.600 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.610 1496.000 1454.890 1500.000 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1374.320 4.000 1374.920 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1391.320 4.000 1391.920 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1474.960 1500.000 1475.560 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.550 1496.000 1472.830 1500.000 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.470 0.000 1473.750 4.000 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1440.960 4.000 1441.560 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 1496.000 1490.770 1500.000 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.280 4.000 1491.880 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 1496.000 352.270 1500.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 414.840 1500.000 415.440 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 496.440 1500.000 497.040 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 1496.000 478.770 1500.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 529.080 1500.000 529.680 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 1496.000 568.930 1500.000 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 610.680 1500.000 611.280 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 1496.000 605.270 1500.000 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 675.960 1500.000 676.560 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 692.280 1500.000 692.880 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.280 4.000 641.880 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 1496.000 623.210 1500.000 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 1496.000 641.610 1500.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 1496.000 659.550 1500.000 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 0.000 803.070 4.000 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 0.000 820.550 4.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 773.200 1500.000 773.800 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 805.840 1500.000 806.440 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 822.160 1500.000 822.760 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 838.480 1500.000 839.080 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 854.800 1500.000 855.400 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 1496.000 768.110 1500.000 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 1496.000 153.550 1500.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 791.560 4.000 792.160 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 871.120 1500.000 871.720 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 1496.000 840.330 1500.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.200 4.000 841.800 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 903.760 1500.000 904.360 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 1496.000 858.270 1500.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 4.000 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 0.000 961.770 4.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 0.000 997.190 4.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 153.720 1500.000 154.320 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 874.520 4.000 875.120 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 891.520 4.000 892.120 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 1496.000 930.490 1500.000 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 0.000 1032.610 4.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 1496.000 966.830 1500.000 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 4.000 975.080 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 991.480 4.000 992.080 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 0.000 1067.570 4.000 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 1496.000 1002.710 1500.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1018.000 1500.000 1018.600 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 0.000 1102.990 4.000 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.120 4.000 1041.720 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 1496.000 1021.110 1500.000 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 1496.000 1056.990 1500.000 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1034.320 1500.000 1034.920 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1066.960 1500.000 1067.560 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1058.120 4.000 1058.720 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1107.760 4.000 1108.360 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.610 0.000 1155.890 4.000 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.760 4.000 1125.360 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1099.600 1500.000 1100.200 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.080 4.000 1141.680 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1132.240 1500.000 1132.840 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1148.560 1500.000 1149.160 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1164.880 1500.000 1165.480 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 1496.000 262.110 1500.000 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1197.520 1500.000 1198.120 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1230.160 1500.000 1230.760 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1246.480 1500.000 1247.080 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1262.800 1500.000 1263.400 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1174.400 4.000 1175.000 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1191.400 4.000 1192.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.720 4.000 1208.320 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.450 0.000 1226.730 4.000 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.610 1496.000 1201.890 1500.000 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 235.320 1500.000 235.920 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 1496.000 9.110 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 1496.000 27.050 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 39.480 1500.000 40.080 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 1496.000 297.990 1500.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 284.280 1500.000 284.880 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 300.600 1500.000 301.200 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 365.880 1500.000 366.480 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 431.160 1500.000 431.760 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 1496.000 424.490 1500.000 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 1496.000 442.430 1500.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 512.760 1500.000 513.360 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 1496.000 533.050 1500.000 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 578.040 1500.000 578.640 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 627.000 1500.000 627.600 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 659.640 1500.000 660.240 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 1496.000 117.210 1500.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 708.600 1500.000 709.200 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1496.000 135.610 1500.000 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 121.080 1500.000 121.680 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 1496.000 189.430 1500.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 1496.000 243.710 1500.000 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 4.000 325.000 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1494.855 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.915 1488.080 ;
      LAYER met2 ;
        RECT 6.990 1495.720 8.550 1496.410 ;
        RECT 9.390 1495.720 26.490 1496.410 ;
        RECT 27.330 1495.720 44.430 1496.410 ;
        RECT 45.270 1495.720 62.370 1496.410 ;
        RECT 63.210 1495.720 80.770 1496.410 ;
        RECT 81.610 1495.720 98.710 1496.410 ;
        RECT 99.550 1495.720 116.650 1496.410 ;
        RECT 117.490 1495.720 135.050 1496.410 ;
        RECT 135.890 1495.720 152.990 1496.410 ;
        RECT 153.830 1495.720 170.930 1496.410 ;
        RECT 171.770 1495.720 188.870 1496.410 ;
        RECT 189.710 1495.720 207.270 1496.410 ;
        RECT 208.110 1495.720 225.210 1496.410 ;
        RECT 226.050 1495.720 243.150 1496.410 ;
        RECT 243.990 1495.720 261.550 1496.410 ;
        RECT 262.390 1495.720 279.490 1496.410 ;
        RECT 280.330 1495.720 297.430 1496.410 ;
        RECT 298.270 1495.720 315.370 1496.410 ;
        RECT 316.210 1495.720 333.770 1496.410 ;
        RECT 334.610 1495.720 351.710 1496.410 ;
        RECT 352.550 1495.720 369.650 1496.410 ;
        RECT 370.490 1495.720 388.050 1496.410 ;
        RECT 388.890 1495.720 405.990 1496.410 ;
        RECT 406.830 1495.720 423.930 1496.410 ;
        RECT 424.770 1495.720 441.870 1496.410 ;
        RECT 442.710 1495.720 460.270 1496.410 ;
        RECT 461.110 1495.720 478.210 1496.410 ;
        RECT 479.050 1495.720 496.150 1496.410 ;
        RECT 496.990 1495.720 514.550 1496.410 ;
        RECT 515.390 1495.720 532.490 1496.410 ;
        RECT 533.330 1495.720 550.430 1496.410 ;
        RECT 551.270 1495.720 568.370 1496.410 ;
        RECT 569.210 1495.720 586.770 1496.410 ;
        RECT 587.610 1495.720 604.710 1496.410 ;
        RECT 605.550 1495.720 622.650 1496.410 ;
        RECT 623.490 1495.720 641.050 1496.410 ;
        RECT 641.890 1495.720 658.990 1496.410 ;
        RECT 659.830 1495.720 676.930 1496.410 ;
        RECT 677.770 1495.720 694.870 1496.410 ;
        RECT 695.710 1495.720 713.270 1496.410 ;
        RECT 714.110 1495.720 731.210 1496.410 ;
        RECT 732.050 1495.720 749.150 1496.410 ;
        RECT 749.990 1495.720 767.550 1496.410 ;
        RECT 768.390 1495.720 785.490 1496.410 ;
        RECT 786.330 1495.720 803.430 1496.410 ;
        RECT 804.270 1495.720 821.830 1496.410 ;
        RECT 822.670 1495.720 839.770 1496.410 ;
        RECT 840.610 1495.720 857.710 1496.410 ;
        RECT 858.550 1495.720 875.650 1496.410 ;
        RECT 876.490 1495.720 894.050 1496.410 ;
        RECT 894.890 1495.720 911.990 1496.410 ;
        RECT 912.830 1495.720 929.930 1496.410 ;
        RECT 930.770 1495.720 948.330 1496.410 ;
        RECT 949.170 1495.720 966.270 1496.410 ;
        RECT 967.110 1495.720 984.210 1496.410 ;
        RECT 985.050 1495.720 1002.150 1496.410 ;
        RECT 1002.990 1495.720 1020.550 1496.410 ;
        RECT 1021.390 1495.720 1038.490 1496.410 ;
        RECT 1039.330 1495.720 1056.430 1496.410 ;
        RECT 1057.270 1495.720 1074.830 1496.410 ;
        RECT 1075.670 1495.720 1092.770 1496.410 ;
        RECT 1093.610 1495.720 1110.710 1496.410 ;
        RECT 1111.550 1495.720 1128.650 1496.410 ;
        RECT 1129.490 1495.720 1147.050 1496.410 ;
        RECT 1147.890 1495.720 1164.990 1496.410 ;
        RECT 1165.830 1495.720 1182.930 1496.410 ;
        RECT 1183.770 1495.720 1201.330 1496.410 ;
        RECT 1202.170 1495.720 1219.270 1496.410 ;
        RECT 1220.110 1495.720 1237.210 1496.410 ;
        RECT 1238.050 1495.720 1255.150 1496.410 ;
        RECT 1255.990 1495.720 1273.550 1496.410 ;
        RECT 1274.390 1495.720 1291.490 1496.410 ;
        RECT 1292.330 1495.720 1309.430 1496.410 ;
        RECT 1310.270 1495.720 1327.830 1496.410 ;
        RECT 1328.670 1495.720 1345.770 1496.410 ;
        RECT 1346.610 1495.720 1363.710 1496.410 ;
        RECT 1364.550 1495.720 1381.650 1496.410 ;
        RECT 1382.490 1495.720 1400.050 1496.410 ;
        RECT 1400.890 1495.720 1417.990 1496.410 ;
        RECT 1418.830 1495.720 1435.930 1496.410 ;
        RECT 1436.770 1495.720 1454.330 1496.410 ;
        RECT 1455.170 1495.720 1472.270 1496.410 ;
        RECT 1473.110 1495.720 1490.210 1496.410 ;
        RECT 1491.050 1495.720 1491.220 1496.410 ;
        RECT 6.990 4.280 1491.220 1495.720 ;
        RECT 6.990 3.670 8.550 4.280 ;
        RECT 9.390 3.670 26.030 4.280 ;
        RECT 26.870 3.670 43.510 4.280 ;
        RECT 44.350 3.670 61.450 4.280 ;
        RECT 62.290 3.670 78.930 4.280 ;
        RECT 79.770 3.670 96.410 4.280 ;
        RECT 97.250 3.670 114.350 4.280 ;
        RECT 115.190 3.670 131.830 4.280 ;
        RECT 132.670 3.670 149.310 4.280 ;
        RECT 150.150 3.670 167.250 4.280 ;
        RECT 168.090 3.670 184.730 4.280 ;
        RECT 185.570 3.670 202.670 4.280 ;
        RECT 203.510 3.670 220.150 4.280 ;
        RECT 220.990 3.670 237.630 4.280 ;
        RECT 238.470 3.670 255.570 4.280 ;
        RECT 256.410 3.670 273.050 4.280 ;
        RECT 273.890 3.670 290.530 4.280 ;
        RECT 291.370 3.670 308.470 4.280 ;
        RECT 309.310 3.670 325.950 4.280 ;
        RECT 326.790 3.670 343.430 4.280 ;
        RECT 344.270 3.670 361.370 4.280 ;
        RECT 362.210 3.670 378.850 4.280 ;
        RECT 379.690 3.670 396.790 4.280 ;
        RECT 397.630 3.670 414.270 4.280 ;
        RECT 415.110 3.670 431.750 4.280 ;
        RECT 432.590 3.670 449.690 4.280 ;
        RECT 450.530 3.670 467.170 4.280 ;
        RECT 468.010 3.670 484.650 4.280 ;
        RECT 485.490 3.670 502.590 4.280 ;
        RECT 503.430 3.670 520.070 4.280 ;
        RECT 520.910 3.670 537.550 4.280 ;
        RECT 538.390 3.670 555.490 4.280 ;
        RECT 556.330 3.670 572.970 4.280 ;
        RECT 573.810 3.670 590.910 4.280 ;
        RECT 591.750 3.670 608.390 4.280 ;
        RECT 609.230 3.670 625.870 4.280 ;
        RECT 626.710 3.670 643.810 4.280 ;
        RECT 644.650 3.670 661.290 4.280 ;
        RECT 662.130 3.670 678.770 4.280 ;
        RECT 679.610 3.670 696.710 4.280 ;
        RECT 697.550 3.670 714.190 4.280 ;
        RECT 715.030 3.670 731.670 4.280 ;
        RECT 732.510 3.670 749.610 4.280 ;
        RECT 750.450 3.670 767.090 4.280 ;
        RECT 767.930 3.670 785.030 4.280 ;
        RECT 785.870 3.670 802.510 4.280 ;
        RECT 803.350 3.670 819.990 4.280 ;
        RECT 820.830 3.670 837.930 4.280 ;
        RECT 838.770 3.670 855.410 4.280 ;
        RECT 856.250 3.670 872.890 4.280 ;
        RECT 873.730 3.670 890.830 4.280 ;
        RECT 891.670 3.670 908.310 4.280 ;
        RECT 909.150 3.670 925.790 4.280 ;
        RECT 926.630 3.670 943.730 4.280 ;
        RECT 944.570 3.670 961.210 4.280 ;
        RECT 962.050 3.670 979.150 4.280 ;
        RECT 979.990 3.670 996.630 4.280 ;
        RECT 997.470 3.670 1014.110 4.280 ;
        RECT 1014.950 3.670 1032.050 4.280 ;
        RECT 1032.890 3.670 1049.530 4.280 ;
        RECT 1050.370 3.670 1067.010 4.280 ;
        RECT 1067.850 3.670 1084.950 4.280 ;
        RECT 1085.790 3.670 1102.430 4.280 ;
        RECT 1103.270 3.670 1119.910 4.280 ;
        RECT 1120.750 3.670 1137.850 4.280 ;
        RECT 1138.690 3.670 1155.330 4.280 ;
        RECT 1156.170 3.670 1173.270 4.280 ;
        RECT 1174.110 3.670 1190.750 4.280 ;
        RECT 1191.590 3.670 1208.230 4.280 ;
        RECT 1209.070 3.670 1226.170 4.280 ;
        RECT 1227.010 3.670 1243.650 4.280 ;
        RECT 1244.490 3.670 1261.130 4.280 ;
        RECT 1261.970 3.670 1279.070 4.280 ;
        RECT 1279.910 3.670 1296.550 4.280 ;
        RECT 1297.390 3.670 1314.030 4.280 ;
        RECT 1314.870 3.670 1331.970 4.280 ;
        RECT 1332.810 3.670 1349.450 4.280 ;
        RECT 1350.290 3.670 1367.390 4.280 ;
        RECT 1368.230 3.670 1384.870 4.280 ;
        RECT 1385.710 3.670 1402.350 4.280 ;
        RECT 1403.190 3.670 1420.290 4.280 ;
        RECT 1421.130 3.670 1437.770 4.280 ;
        RECT 1438.610 3.670 1455.250 4.280 ;
        RECT 1456.090 3.670 1473.190 4.280 ;
        RECT 1474.030 3.670 1490.670 4.280 ;
      LAYER met3 ;
        RECT 4.400 1490.880 1495.600 1491.745 ;
        RECT 4.000 1475.960 1496.000 1490.880 ;
        RECT 4.000 1475.280 1495.600 1475.960 ;
        RECT 4.400 1474.560 1495.600 1475.280 ;
        RECT 4.400 1473.880 1496.000 1474.560 ;
        RECT 4.000 1459.640 1496.000 1473.880 ;
        RECT 4.000 1458.960 1495.600 1459.640 ;
        RECT 4.400 1458.240 1495.600 1458.960 ;
        RECT 4.400 1457.560 1496.000 1458.240 ;
        RECT 4.000 1443.320 1496.000 1457.560 ;
        RECT 4.000 1441.960 1495.600 1443.320 ;
        RECT 4.400 1441.920 1495.600 1441.960 ;
        RECT 4.400 1440.560 1496.000 1441.920 ;
        RECT 4.000 1427.000 1496.000 1440.560 ;
        RECT 4.000 1425.640 1495.600 1427.000 ;
        RECT 4.400 1425.600 1495.600 1425.640 ;
        RECT 4.400 1424.240 1496.000 1425.600 ;
        RECT 4.000 1410.680 1496.000 1424.240 ;
        RECT 4.000 1409.280 1495.600 1410.680 ;
        RECT 4.000 1408.640 1496.000 1409.280 ;
        RECT 4.400 1407.240 1496.000 1408.640 ;
        RECT 4.000 1394.360 1496.000 1407.240 ;
        RECT 4.000 1392.960 1495.600 1394.360 ;
        RECT 4.000 1392.320 1496.000 1392.960 ;
        RECT 4.400 1390.920 1496.000 1392.320 ;
        RECT 4.000 1378.040 1496.000 1390.920 ;
        RECT 4.000 1376.640 1495.600 1378.040 ;
        RECT 4.000 1375.320 1496.000 1376.640 ;
        RECT 4.400 1373.920 1496.000 1375.320 ;
        RECT 4.000 1361.720 1496.000 1373.920 ;
        RECT 4.000 1360.320 1495.600 1361.720 ;
        RECT 4.000 1359.000 1496.000 1360.320 ;
        RECT 4.400 1357.600 1496.000 1359.000 ;
        RECT 4.000 1345.400 1496.000 1357.600 ;
        RECT 4.000 1344.000 1495.600 1345.400 ;
        RECT 4.000 1342.000 1496.000 1344.000 ;
        RECT 4.400 1340.600 1496.000 1342.000 ;
        RECT 4.000 1329.080 1496.000 1340.600 ;
        RECT 4.000 1327.680 1495.600 1329.080 ;
        RECT 4.000 1325.680 1496.000 1327.680 ;
        RECT 4.400 1324.280 1496.000 1325.680 ;
        RECT 4.000 1312.760 1496.000 1324.280 ;
        RECT 4.000 1311.360 1495.600 1312.760 ;
        RECT 4.000 1308.680 1496.000 1311.360 ;
        RECT 4.400 1307.280 1496.000 1308.680 ;
        RECT 4.000 1296.440 1496.000 1307.280 ;
        RECT 4.000 1295.040 1495.600 1296.440 ;
        RECT 4.000 1292.360 1496.000 1295.040 ;
        RECT 4.400 1290.960 1496.000 1292.360 ;
        RECT 4.000 1280.120 1496.000 1290.960 ;
        RECT 4.000 1278.720 1495.600 1280.120 ;
        RECT 4.000 1275.360 1496.000 1278.720 ;
        RECT 4.400 1273.960 1496.000 1275.360 ;
        RECT 4.000 1263.800 1496.000 1273.960 ;
        RECT 4.000 1262.400 1495.600 1263.800 ;
        RECT 4.000 1259.040 1496.000 1262.400 ;
        RECT 4.400 1257.640 1496.000 1259.040 ;
        RECT 4.000 1247.480 1496.000 1257.640 ;
        RECT 4.000 1246.080 1495.600 1247.480 ;
        RECT 4.000 1242.040 1496.000 1246.080 ;
        RECT 4.400 1240.640 1496.000 1242.040 ;
        RECT 4.000 1231.160 1496.000 1240.640 ;
        RECT 4.000 1229.760 1495.600 1231.160 ;
        RECT 4.000 1225.720 1496.000 1229.760 ;
        RECT 4.400 1224.320 1496.000 1225.720 ;
        RECT 4.000 1214.840 1496.000 1224.320 ;
        RECT 4.000 1213.440 1495.600 1214.840 ;
        RECT 4.000 1208.720 1496.000 1213.440 ;
        RECT 4.400 1207.320 1496.000 1208.720 ;
        RECT 4.000 1198.520 1496.000 1207.320 ;
        RECT 4.000 1197.120 1495.600 1198.520 ;
        RECT 4.000 1192.400 1496.000 1197.120 ;
        RECT 4.400 1191.000 1496.000 1192.400 ;
        RECT 4.000 1182.200 1496.000 1191.000 ;
        RECT 4.000 1180.800 1495.600 1182.200 ;
        RECT 4.000 1175.400 1496.000 1180.800 ;
        RECT 4.400 1174.000 1496.000 1175.400 ;
        RECT 4.000 1165.880 1496.000 1174.000 ;
        RECT 4.000 1164.480 1495.600 1165.880 ;
        RECT 4.000 1159.080 1496.000 1164.480 ;
        RECT 4.400 1157.680 1496.000 1159.080 ;
        RECT 4.000 1149.560 1496.000 1157.680 ;
        RECT 4.000 1148.160 1495.600 1149.560 ;
        RECT 4.000 1142.080 1496.000 1148.160 ;
        RECT 4.400 1140.680 1496.000 1142.080 ;
        RECT 4.000 1133.240 1496.000 1140.680 ;
        RECT 4.000 1131.840 1495.600 1133.240 ;
        RECT 4.000 1125.760 1496.000 1131.840 ;
        RECT 4.400 1124.360 1496.000 1125.760 ;
        RECT 4.000 1116.920 1496.000 1124.360 ;
        RECT 4.000 1115.520 1495.600 1116.920 ;
        RECT 4.000 1108.760 1496.000 1115.520 ;
        RECT 4.400 1107.360 1496.000 1108.760 ;
        RECT 4.000 1100.600 1496.000 1107.360 ;
        RECT 4.000 1099.200 1495.600 1100.600 ;
        RECT 4.000 1092.440 1496.000 1099.200 ;
        RECT 4.400 1091.040 1496.000 1092.440 ;
        RECT 4.000 1084.280 1496.000 1091.040 ;
        RECT 4.000 1082.880 1495.600 1084.280 ;
        RECT 4.000 1075.440 1496.000 1082.880 ;
        RECT 4.400 1074.040 1496.000 1075.440 ;
        RECT 4.000 1067.960 1496.000 1074.040 ;
        RECT 4.000 1066.560 1495.600 1067.960 ;
        RECT 4.000 1059.120 1496.000 1066.560 ;
        RECT 4.400 1057.720 1496.000 1059.120 ;
        RECT 4.000 1051.640 1496.000 1057.720 ;
        RECT 4.000 1050.240 1495.600 1051.640 ;
        RECT 4.000 1042.120 1496.000 1050.240 ;
        RECT 4.400 1040.720 1496.000 1042.120 ;
        RECT 4.000 1035.320 1496.000 1040.720 ;
        RECT 4.000 1033.920 1495.600 1035.320 ;
        RECT 4.000 1025.800 1496.000 1033.920 ;
        RECT 4.400 1024.400 1496.000 1025.800 ;
        RECT 4.000 1019.000 1496.000 1024.400 ;
        RECT 4.000 1017.600 1495.600 1019.000 ;
        RECT 4.000 1008.800 1496.000 1017.600 ;
        RECT 4.400 1007.400 1496.000 1008.800 ;
        RECT 4.000 1002.680 1496.000 1007.400 ;
        RECT 4.000 1001.280 1495.600 1002.680 ;
        RECT 4.000 992.480 1496.000 1001.280 ;
        RECT 4.400 991.080 1496.000 992.480 ;
        RECT 4.000 986.360 1496.000 991.080 ;
        RECT 4.000 984.960 1495.600 986.360 ;
        RECT 4.000 975.480 1496.000 984.960 ;
        RECT 4.400 974.080 1496.000 975.480 ;
        RECT 4.000 970.040 1496.000 974.080 ;
        RECT 4.000 968.640 1495.600 970.040 ;
        RECT 4.000 959.160 1496.000 968.640 ;
        RECT 4.400 957.760 1496.000 959.160 ;
        RECT 4.000 953.720 1496.000 957.760 ;
        RECT 4.000 952.320 1495.600 953.720 ;
        RECT 4.000 942.160 1496.000 952.320 ;
        RECT 4.400 940.760 1496.000 942.160 ;
        RECT 4.000 937.400 1496.000 940.760 ;
        RECT 4.000 936.000 1495.600 937.400 ;
        RECT 4.000 925.840 1496.000 936.000 ;
        RECT 4.400 924.440 1496.000 925.840 ;
        RECT 4.000 921.080 1496.000 924.440 ;
        RECT 4.000 919.680 1495.600 921.080 ;
        RECT 4.000 908.840 1496.000 919.680 ;
        RECT 4.400 907.440 1496.000 908.840 ;
        RECT 4.000 904.760 1496.000 907.440 ;
        RECT 4.000 903.360 1495.600 904.760 ;
        RECT 4.000 892.520 1496.000 903.360 ;
        RECT 4.400 891.120 1496.000 892.520 ;
        RECT 4.000 888.440 1496.000 891.120 ;
        RECT 4.000 887.040 1495.600 888.440 ;
        RECT 4.000 875.520 1496.000 887.040 ;
        RECT 4.400 874.120 1496.000 875.520 ;
        RECT 4.000 872.120 1496.000 874.120 ;
        RECT 4.000 870.720 1495.600 872.120 ;
        RECT 4.000 859.200 1496.000 870.720 ;
        RECT 4.400 857.800 1496.000 859.200 ;
        RECT 4.000 855.800 1496.000 857.800 ;
        RECT 4.000 854.400 1495.600 855.800 ;
        RECT 4.000 842.200 1496.000 854.400 ;
        RECT 4.400 840.800 1496.000 842.200 ;
        RECT 4.000 839.480 1496.000 840.800 ;
        RECT 4.000 838.080 1495.600 839.480 ;
        RECT 4.000 825.880 1496.000 838.080 ;
        RECT 4.400 824.480 1496.000 825.880 ;
        RECT 4.000 823.160 1496.000 824.480 ;
        RECT 4.000 821.760 1495.600 823.160 ;
        RECT 4.000 808.880 1496.000 821.760 ;
        RECT 4.400 807.480 1496.000 808.880 ;
        RECT 4.000 806.840 1496.000 807.480 ;
        RECT 4.000 805.440 1495.600 806.840 ;
        RECT 4.000 792.560 1496.000 805.440 ;
        RECT 4.400 791.160 1496.000 792.560 ;
        RECT 4.000 790.520 1496.000 791.160 ;
        RECT 4.000 789.120 1495.600 790.520 ;
        RECT 4.000 775.560 1496.000 789.120 ;
        RECT 4.400 774.200 1496.000 775.560 ;
        RECT 4.400 774.160 1495.600 774.200 ;
        RECT 4.000 772.800 1495.600 774.160 ;
        RECT 4.000 759.240 1496.000 772.800 ;
        RECT 4.400 758.560 1496.000 759.240 ;
        RECT 4.400 757.840 1495.600 758.560 ;
        RECT 4.000 757.160 1495.600 757.840 ;
        RECT 4.000 742.240 1496.000 757.160 ;
        RECT 4.400 740.840 1495.600 742.240 ;
        RECT 4.000 725.920 1496.000 740.840 ;
        RECT 4.000 725.240 1495.600 725.920 ;
        RECT 4.400 724.520 1495.600 725.240 ;
        RECT 4.400 723.840 1496.000 724.520 ;
        RECT 4.000 709.600 1496.000 723.840 ;
        RECT 4.000 708.920 1495.600 709.600 ;
        RECT 4.400 708.200 1495.600 708.920 ;
        RECT 4.400 707.520 1496.000 708.200 ;
        RECT 4.000 693.280 1496.000 707.520 ;
        RECT 4.000 691.920 1495.600 693.280 ;
        RECT 4.400 691.880 1495.600 691.920 ;
        RECT 4.400 690.520 1496.000 691.880 ;
        RECT 4.000 676.960 1496.000 690.520 ;
        RECT 4.000 675.600 1495.600 676.960 ;
        RECT 4.400 675.560 1495.600 675.600 ;
        RECT 4.400 674.200 1496.000 675.560 ;
        RECT 4.000 660.640 1496.000 674.200 ;
        RECT 4.000 659.240 1495.600 660.640 ;
        RECT 4.000 658.600 1496.000 659.240 ;
        RECT 4.400 657.200 1496.000 658.600 ;
        RECT 4.000 644.320 1496.000 657.200 ;
        RECT 4.000 642.920 1495.600 644.320 ;
        RECT 4.000 642.280 1496.000 642.920 ;
        RECT 4.400 640.880 1496.000 642.280 ;
        RECT 4.000 628.000 1496.000 640.880 ;
        RECT 4.000 626.600 1495.600 628.000 ;
        RECT 4.000 625.280 1496.000 626.600 ;
        RECT 4.400 623.880 1496.000 625.280 ;
        RECT 4.000 611.680 1496.000 623.880 ;
        RECT 4.000 610.280 1495.600 611.680 ;
        RECT 4.000 608.960 1496.000 610.280 ;
        RECT 4.400 607.560 1496.000 608.960 ;
        RECT 4.000 595.360 1496.000 607.560 ;
        RECT 4.000 593.960 1495.600 595.360 ;
        RECT 4.000 591.960 1496.000 593.960 ;
        RECT 4.400 590.560 1496.000 591.960 ;
        RECT 4.000 579.040 1496.000 590.560 ;
        RECT 4.000 577.640 1495.600 579.040 ;
        RECT 4.000 575.640 1496.000 577.640 ;
        RECT 4.400 574.240 1496.000 575.640 ;
        RECT 4.000 562.720 1496.000 574.240 ;
        RECT 4.000 561.320 1495.600 562.720 ;
        RECT 4.000 558.640 1496.000 561.320 ;
        RECT 4.400 557.240 1496.000 558.640 ;
        RECT 4.000 546.400 1496.000 557.240 ;
        RECT 4.000 545.000 1495.600 546.400 ;
        RECT 4.000 542.320 1496.000 545.000 ;
        RECT 4.400 540.920 1496.000 542.320 ;
        RECT 4.000 530.080 1496.000 540.920 ;
        RECT 4.000 528.680 1495.600 530.080 ;
        RECT 4.000 525.320 1496.000 528.680 ;
        RECT 4.400 523.920 1496.000 525.320 ;
        RECT 4.000 513.760 1496.000 523.920 ;
        RECT 4.000 512.360 1495.600 513.760 ;
        RECT 4.000 509.000 1496.000 512.360 ;
        RECT 4.400 507.600 1496.000 509.000 ;
        RECT 4.000 497.440 1496.000 507.600 ;
        RECT 4.000 496.040 1495.600 497.440 ;
        RECT 4.000 492.000 1496.000 496.040 ;
        RECT 4.400 490.600 1496.000 492.000 ;
        RECT 4.000 481.120 1496.000 490.600 ;
        RECT 4.000 479.720 1495.600 481.120 ;
        RECT 4.000 475.680 1496.000 479.720 ;
        RECT 4.400 474.280 1496.000 475.680 ;
        RECT 4.000 464.800 1496.000 474.280 ;
        RECT 4.000 463.400 1495.600 464.800 ;
        RECT 4.000 458.680 1496.000 463.400 ;
        RECT 4.400 457.280 1496.000 458.680 ;
        RECT 4.000 448.480 1496.000 457.280 ;
        RECT 4.000 447.080 1495.600 448.480 ;
        RECT 4.000 442.360 1496.000 447.080 ;
        RECT 4.400 440.960 1496.000 442.360 ;
        RECT 4.000 432.160 1496.000 440.960 ;
        RECT 4.000 430.760 1495.600 432.160 ;
        RECT 4.000 425.360 1496.000 430.760 ;
        RECT 4.400 423.960 1496.000 425.360 ;
        RECT 4.000 415.840 1496.000 423.960 ;
        RECT 4.000 414.440 1495.600 415.840 ;
        RECT 4.000 409.040 1496.000 414.440 ;
        RECT 4.400 407.640 1496.000 409.040 ;
        RECT 4.000 399.520 1496.000 407.640 ;
        RECT 4.000 398.120 1495.600 399.520 ;
        RECT 4.000 392.040 1496.000 398.120 ;
        RECT 4.400 390.640 1496.000 392.040 ;
        RECT 4.000 383.200 1496.000 390.640 ;
        RECT 4.000 381.800 1495.600 383.200 ;
        RECT 4.000 375.720 1496.000 381.800 ;
        RECT 4.400 374.320 1496.000 375.720 ;
        RECT 4.000 366.880 1496.000 374.320 ;
        RECT 4.000 365.480 1495.600 366.880 ;
        RECT 4.000 358.720 1496.000 365.480 ;
        RECT 4.400 357.320 1496.000 358.720 ;
        RECT 4.000 350.560 1496.000 357.320 ;
        RECT 4.000 349.160 1495.600 350.560 ;
        RECT 4.000 342.400 1496.000 349.160 ;
        RECT 4.400 341.000 1496.000 342.400 ;
        RECT 4.000 334.240 1496.000 341.000 ;
        RECT 4.000 332.840 1495.600 334.240 ;
        RECT 4.000 325.400 1496.000 332.840 ;
        RECT 4.400 324.000 1496.000 325.400 ;
        RECT 4.000 317.920 1496.000 324.000 ;
        RECT 4.000 316.520 1495.600 317.920 ;
        RECT 4.000 309.080 1496.000 316.520 ;
        RECT 4.400 307.680 1496.000 309.080 ;
        RECT 4.000 301.600 1496.000 307.680 ;
        RECT 4.000 300.200 1495.600 301.600 ;
        RECT 4.000 292.080 1496.000 300.200 ;
        RECT 4.400 290.680 1496.000 292.080 ;
        RECT 4.000 285.280 1496.000 290.680 ;
        RECT 4.000 283.880 1495.600 285.280 ;
        RECT 4.000 275.760 1496.000 283.880 ;
        RECT 4.400 274.360 1496.000 275.760 ;
        RECT 4.000 268.960 1496.000 274.360 ;
        RECT 4.000 267.560 1495.600 268.960 ;
        RECT 4.000 258.760 1496.000 267.560 ;
        RECT 4.400 257.360 1496.000 258.760 ;
        RECT 4.000 252.640 1496.000 257.360 ;
        RECT 4.000 251.240 1495.600 252.640 ;
        RECT 4.000 242.440 1496.000 251.240 ;
        RECT 4.400 241.040 1496.000 242.440 ;
        RECT 4.000 236.320 1496.000 241.040 ;
        RECT 4.000 234.920 1495.600 236.320 ;
        RECT 4.000 225.440 1496.000 234.920 ;
        RECT 4.400 224.040 1496.000 225.440 ;
        RECT 4.000 220.000 1496.000 224.040 ;
        RECT 4.000 218.600 1495.600 220.000 ;
        RECT 4.000 209.120 1496.000 218.600 ;
        RECT 4.400 207.720 1496.000 209.120 ;
        RECT 4.000 203.680 1496.000 207.720 ;
        RECT 4.000 202.280 1495.600 203.680 ;
        RECT 4.000 192.120 1496.000 202.280 ;
        RECT 4.400 190.720 1496.000 192.120 ;
        RECT 4.000 187.360 1496.000 190.720 ;
        RECT 4.000 185.960 1495.600 187.360 ;
        RECT 4.000 175.800 1496.000 185.960 ;
        RECT 4.400 174.400 1496.000 175.800 ;
        RECT 4.000 171.040 1496.000 174.400 ;
        RECT 4.000 169.640 1495.600 171.040 ;
        RECT 4.000 158.800 1496.000 169.640 ;
        RECT 4.400 157.400 1496.000 158.800 ;
        RECT 4.000 154.720 1496.000 157.400 ;
        RECT 4.000 153.320 1495.600 154.720 ;
        RECT 4.000 142.480 1496.000 153.320 ;
        RECT 4.400 141.080 1496.000 142.480 ;
        RECT 4.000 138.400 1496.000 141.080 ;
        RECT 4.000 137.000 1495.600 138.400 ;
        RECT 4.000 125.480 1496.000 137.000 ;
        RECT 4.400 124.080 1496.000 125.480 ;
        RECT 4.000 122.080 1496.000 124.080 ;
        RECT 4.000 120.680 1495.600 122.080 ;
        RECT 4.000 109.160 1496.000 120.680 ;
        RECT 4.400 107.760 1496.000 109.160 ;
        RECT 4.000 105.760 1496.000 107.760 ;
        RECT 4.000 104.360 1495.600 105.760 ;
        RECT 4.000 92.160 1496.000 104.360 ;
        RECT 4.400 90.760 1496.000 92.160 ;
        RECT 4.000 89.440 1496.000 90.760 ;
        RECT 4.000 88.040 1495.600 89.440 ;
        RECT 4.000 75.840 1496.000 88.040 ;
        RECT 4.400 74.440 1496.000 75.840 ;
        RECT 4.000 73.120 1496.000 74.440 ;
        RECT 4.000 71.720 1495.600 73.120 ;
        RECT 4.000 58.840 1496.000 71.720 ;
        RECT 4.400 57.440 1496.000 58.840 ;
        RECT 4.000 56.800 1496.000 57.440 ;
        RECT 4.000 55.400 1495.600 56.800 ;
        RECT 4.000 42.520 1496.000 55.400 ;
        RECT 4.400 41.120 1496.000 42.520 ;
        RECT 4.000 40.480 1496.000 41.120 ;
        RECT 4.000 39.080 1495.600 40.480 ;
        RECT 4.000 25.520 1496.000 39.080 ;
        RECT 4.400 24.160 1496.000 25.520 ;
        RECT 4.400 24.120 1495.600 24.160 ;
        RECT 4.000 22.760 1495.600 24.120 ;
        RECT 4.000 9.200 1496.000 22.760 ;
        RECT 4.400 8.520 1496.000 9.200 ;
        RECT 4.400 7.800 1495.600 8.520 ;
        RECT 4.000 7.655 1495.600 7.800 ;
      LAYER met4 ;
        RECT 88.615 11.055 97.440 1485.625 ;
        RECT 99.840 11.055 174.240 1485.625 ;
        RECT 176.640 11.055 251.040 1485.625 ;
        RECT 253.440 11.055 327.840 1485.625 ;
        RECT 330.240 11.055 404.640 1485.625 ;
        RECT 407.040 11.055 481.440 1485.625 ;
        RECT 483.840 11.055 558.240 1485.625 ;
        RECT 560.640 11.055 635.040 1485.625 ;
        RECT 637.440 11.055 711.840 1485.625 ;
        RECT 714.240 11.055 788.640 1485.625 ;
        RECT 791.040 11.055 865.440 1485.625 ;
        RECT 867.840 11.055 942.240 1485.625 ;
        RECT 944.640 11.055 1019.040 1485.625 ;
        RECT 1021.440 11.055 1095.840 1485.625 ;
        RECT 1098.240 11.055 1172.640 1485.625 ;
        RECT 1175.040 11.055 1249.440 1485.625 ;
        RECT 1251.840 11.055 1303.345 1485.625 ;
  END
END core
END LIBRARY

