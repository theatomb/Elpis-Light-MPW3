VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.840 4.000 1214.440 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1292.040 1500.000 1292.640 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.710 0.000 1286.990 4.000 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.970 0.000 1324.250 4.000 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1328.080 1500.000 1328.680 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1246.480 4.000 1247.080 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.630 0.000 1379.910 4.000 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1262.800 4.000 1263.400 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1364.120 1500.000 1364.720 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 1496.000 326.970 1500.000 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1400.160 1500.000 1400.760 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.350 1496.000 1348.630 1500.000 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1295.440 4.000 1296.040 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1328.080 4.000 1328.680 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 1496.000 1364.270 1500.000 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 1496.000 1380.370 1500.000 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.430 0.000 1416.710 4.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.830 1496.000 1412.110 1500.000 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.030 1496.000 1444.310 1500.000 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 207.440 1500.000 208.040 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.680 4.000 1410.280 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1442.320 4.000 1442.920 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.670 1496.000 1459.950 1500.000 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1474.960 4.000 1475.560 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 0.000 1453.970 4.000 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.490 0.000 1490.770 4.000 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1472.240 1500.000 1472.840 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.870 1496.000 1492.150 1500.000 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 279.520 1500.000 280.120 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 1496.000 374.810 1500.000 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 1496.000 390.910 1500.000 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 1496.000 454.850 1500.000 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 1496.000 470.950 1500.000 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 8.880 1500.000 9.480 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 1496.000 534.430 1500.000 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 1496.000 582.270 1500.000 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 496.440 1500.000 497.040 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 532.480 1500.000 533.080 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 568.520 1500.000 569.120 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 622.920 1500.000 623.520 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 1496.000 630.110 1500.000 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 677.320 1500.000 677.920 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 713.360 1500.000 713.960 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 1496.000 694.050 1500.000 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 1496.000 726.250 1500.000 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 767.760 1500.000 768.360 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 1496.000 741.890 1500.000 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 803.800 1500.000 804.400 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 822.160 1500.000 822.760 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 1496.000 757.990 1500.000 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 1496.000 774.090 1500.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 0.000 842.630 4.000 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 1496.000 805.830 1500.000 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 875.880 1500.000 876.480 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 894.240 1500.000 894.840 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 1496.000 837.570 1500.000 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 948.640 1500.000 949.240 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 966.320 1500.000 966.920 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 1496.000 869.770 1500.000 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1002.360 1500.000 1002.960 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 1496.000 885.870 1500.000 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 789.520 4.000 790.120 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 1496.000 231.290 1500.000 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 1496.000 901.510 1500.000 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.070 0.000 972.350 4.000 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 1496.000 933.710 1500.000 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1056.760 1500.000 1057.360 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 1496.000 949.350 1500.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 0.000 990.750 4.000 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 0.000 1009.610 4.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 838.480 4.000 839.080 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.730 0.000 1028.010 4.000 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 98.640 1500.000 99.240 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.390 0.000 1083.670 4.000 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 1496.000 997.190 1500.000 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 1496.000 1029.390 1500.000 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 0.000 1102.070 4.000 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 1496.000 1045.030 1500.000 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1128.840 1500.000 1129.440 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.590 0.000 1138.870 4.000 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1147.200 1500.000 1147.800 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.450 0.000 1157.730 4.000 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 1496.000 1077.230 1500.000 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.050 1496.000 1093.330 1500.000 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.000 4.000 1018.600 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.960 4.000 1067.560 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 1496.000 1125.070 1500.000 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.890 1496.000 1141.170 1500.000 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1165.560 1500.000 1166.160 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1183.240 1500.000 1183.840 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 1496.000 295.230 1500.000 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 1496.000 1172.910 1500.000 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.920 4.000 1116.520 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1219.280 1500.000 1219.880 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1148.560 4.000 1149.160 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1164.880 4.000 1165.480 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 1496.000 1236.850 1500.000 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1181.200 4.000 1181.800 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.310 1496.000 1268.590 1500.000 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1255.320 1500.000 1255.920 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.410 1496.000 1284.690 1500.000 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 1496.000 135.610 1500.000 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 225.120 1500.000 225.720 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 1496.000 359.170 1500.000 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 1496.000 407.010 1500.000 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 315.560 1500.000 316.160 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 1496.000 438.750 1500.000 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 424.360 1500.000 424.960 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 1496.000 167.350 1500.000 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 460.400 1500.000 461.000 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 0.000 602.050 4.000 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 1496.000 614.470 1500.000 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 586.880 1500.000 587.480 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 641.280 1500.000 641.880 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 0.000 676.110 4.000 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 1496.000 678.410 1500.000 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 62.600 1500.000 63.200 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 80.960 1500.000 81.560 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 171.400 1500.000 172.000 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 1496.000 39.930 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 1496.000 87.770 1500.000 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 1496.000 71.670 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 1496.000 103.870 1500.000 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1496.000 119.510 1500.000 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 1496.000 56.030 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 1496.000 151.710 1500.000 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 333.920 1500.000 334.520 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 351.600 1500.000 352.200 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 26.560 1500.000 27.160 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 44.920 1500.000 45.520 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 1496.000 199.550 1500.000 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 1496.000 247.390 1500.000 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 117.000 1500.000 117.600 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 153.040 1500.000 153.640 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.160 4.000 1230.760 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.310 0.000 1268.590 4.000 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.570 0.000 1305.850 4.000 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1300.510 1496.000 1300.790 1500.000 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1309.720 1500.000 1310.320 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 1496.000 1316.430 1500.000 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 0.000 1361.050 4.000 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1345.760 1500.000 1346.360 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.250 1496.000 1332.530 1500.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1381.800 1500.000 1382.400 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.120 4.000 1279.720 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.030 0.000 1398.310 4.000 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1311.760 4.000 1312.360 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1344.400 4.000 1345.000 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1418.520 1500.000 1419.120 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.190 1496.000 1396.470 1500.000 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.720 4.000 1361.320 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1393.360 4.000 1393.960 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.930 1496.000 1428.210 1500.000 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1436.200 1500.000 1436.800 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 243.480 1500.000 244.080 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1426.000 4.000 1426.600 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.830 0.000 1435.110 4.000 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1458.640 4.000 1459.240 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.770 1496.000 1476.050 1500.000 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.090 0.000 1472.370 4.000 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1454.560 1500.000 1455.160 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.280 4.000 1491.880 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1490.600 1500.000 1491.200 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 369.960 1500.000 370.560 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 388.320 1500.000 388.920 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 406.000 1500.000 406.600 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 442.040 1500.000 442.640 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 1496.000 502.690 1500.000 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 1496.000 550.530 1500.000 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 1496.000 598.370 1500.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 605.240 1500.000 605.840 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 658.960 1500.000 659.560 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 1496.000 646.210 1500.000 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 731.720 1500.000 732.320 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 749.400 1500.000 750.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.870 1496.000 710.150 1500.000 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 1496.000 183.450 1500.000 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 785.440 1500.000 786.040 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 0.000 824.230 4.000 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 839.840 1500.000 840.440 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 1496.000 789.730 1500.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 858.200 1500.000 858.800 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.650 1496.000 821.930 1500.000 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.280 4.000 692.880 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 911.920 1500.000 912.520 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 930.280 1500.000 930.880 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 1496.000 853.670 1500.000 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 984.680 1500.000 985.280 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 0.000 898.290 4.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 4.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1020.720 1500.000 1021.320 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 4.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 0.000 953.950 4.000 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 1496.000 263.490 1500.000 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.330 1496.000 917.610 1500.000 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1038.400 1500.000 1039.000 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1075.120 1500.000 1075.720 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.170 1496.000 965.450 1500.000 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.160 4.000 822.760 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 1496.000 981.550 1500.000 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1092.800 1500.000 1093.400 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.800 4.000 855.400 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 135.360 1500.000 135.960 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.120 4.000 871.720 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1111.160 1500.000 1111.760 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 1496.000 1013.290 1500.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.760 4.000 904.360 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 936.400 4.000 937.000 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.720 4.000 953.320 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.850 1496.000 1061.130 1500.000 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 985.360 4.000 985.960 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.680 4.000 1002.280 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1034.320 4.000 1034.920 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.690 1496.000 1108.970 1500.000 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 0.000 1176.130 4.000 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1083.280 4.000 1083.880 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1212.650 0.000 1212.930 4.000 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.530 1496.000 1156.810 1500.000 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1201.600 1500.000 1202.200 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 1496.000 311.330 1500.000 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.730 1496.000 1189.010 1500.000 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1237.640 1500.000 1238.240 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 1496.000 1204.650 1500.000 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 1496.000 1220.750 1500.000 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.510 0.000 1231.790 4.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.210 1496.000 1252.490 1500.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 0.000 1250.190 4.000 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1197.520 4.000 1198.120 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1273.680 1500.000 1274.280 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 1496.000 8.190 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 1496.000 23.830 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 1496.000 343.070 1500.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 261.840 1500.000 262.440 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 297.880 1500.000 298.480 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 1496.000 422.650 1500.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 1496.000 486.590 1500.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 1496.000 518.790 1500.000 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 478.760 1500.000 479.360 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 1496.000 566.630 1500.000 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 514.800 1500.000 515.400 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 550.840 1500.000 551.440 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 1496.000 662.310 1500.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 0.000 712.910 4.000 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 695.000 1500.000 695.600 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 1496.000 215.190 1500.000 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 1496.000 279.130 1500.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 189.080 1500.000 189.680 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.080 1489.160 ;
      LAYER met2 ;
        RECT 6.990 1495.720 7.630 1496.410 ;
        RECT 8.470 1495.720 23.270 1496.410 ;
        RECT 24.110 1495.720 39.370 1496.410 ;
        RECT 40.210 1495.720 55.470 1496.410 ;
        RECT 56.310 1495.720 71.110 1496.410 ;
        RECT 71.950 1495.720 87.210 1496.410 ;
        RECT 88.050 1495.720 103.310 1496.410 ;
        RECT 104.150 1495.720 118.950 1496.410 ;
        RECT 119.790 1495.720 135.050 1496.410 ;
        RECT 135.890 1495.720 151.150 1496.410 ;
        RECT 151.990 1495.720 166.790 1496.410 ;
        RECT 167.630 1495.720 182.890 1496.410 ;
        RECT 183.730 1495.720 198.990 1496.410 ;
        RECT 199.830 1495.720 214.630 1496.410 ;
        RECT 215.470 1495.720 230.730 1496.410 ;
        RECT 231.570 1495.720 246.830 1496.410 ;
        RECT 247.670 1495.720 262.930 1496.410 ;
        RECT 263.770 1495.720 278.570 1496.410 ;
        RECT 279.410 1495.720 294.670 1496.410 ;
        RECT 295.510 1495.720 310.770 1496.410 ;
        RECT 311.610 1495.720 326.410 1496.410 ;
        RECT 327.250 1495.720 342.510 1496.410 ;
        RECT 343.350 1495.720 358.610 1496.410 ;
        RECT 359.450 1495.720 374.250 1496.410 ;
        RECT 375.090 1495.720 390.350 1496.410 ;
        RECT 391.190 1495.720 406.450 1496.410 ;
        RECT 407.290 1495.720 422.090 1496.410 ;
        RECT 422.930 1495.720 438.190 1496.410 ;
        RECT 439.030 1495.720 454.290 1496.410 ;
        RECT 455.130 1495.720 470.390 1496.410 ;
        RECT 471.230 1495.720 486.030 1496.410 ;
        RECT 486.870 1495.720 502.130 1496.410 ;
        RECT 502.970 1495.720 518.230 1496.410 ;
        RECT 519.070 1495.720 533.870 1496.410 ;
        RECT 534.710 1495.720 549.970 1496.410 ;
        RECT 550.810 1495.720 566.070 1496.410 ;
        RECT 566.910 1495.720 581.710 1496.410 ;
        RECT 582.550 1495.720 597.810 1496.410 ;
        RECT 598.650 1495.720 613.910 1496.410 ;
        RECT 614.750 1495.720 629.550 1496.410 ;
        RECT 630.390 1495.720 645.650 1496.410 ;
        RECT 646.490 1495.720 661.750 1496.410 ;
        RECT 662.590 1495.720 677.850 1496.410 ;
        RECT 678.690 1495.720 693.490 1496.410 ;
        RECT 694.330 1495.720 709.590 1496.410 ;
        RECT 710.430 1495.720 725.690 1496.410 ;
        RECT 726.530 1495.720 741.330 1496.410 ;
        RECT 742.170 1495.720 757.430 1496.410 ;
        RECT 758.270 1495.720 773.530 1496.410 ;
        RECT 774.370 1495.720 789.170 1496.410 ;
        RECT 790.010 1495.720 805.270 1496.410 ;
        RECT 806.110 1495.720 821.370 1496.410 ;
        RECT 822.210 1495.720 837.010 1496.410 ;
        RECT 837.850 1495.720 853.110 1496.410 ;
        RECT 853.950 1495.720 869.210 1496.410 ;
        RECT 870.050 1495.720 885.310 1496.410 ;
        RECT 886.150 1495.720 900.950 1496.410 ;
        RECT 901.790 1495.720 917.050 1496.410 ;
        RECT 917.890 1495.720 933.150 1496.410 ;
        RECT 933.990 1495.720 948.790 1496.410 ;
        RECT 949.630 1495.720 964.890 1496.410 ;
        RECT 965.730 1495.720 980.990 1496.410 ;
        RECT 981.830 1495.720 996.630 1496.410 ;
        RECT 997.470 1495.720 1012.730 1496.410 ;
        RECT 1013.570 1495.720 1028.830 1496.410 ;
        RECT 1029.670 1495.720 1044.470 1496.410 ;
        RECT 1045.310 1495.720 1060.570 1496.410 ;
        RECT 1061.410 1495.720 1076.670 1496.410 ;
        RECT 1077.510 1495.720 1092.770 1496.410 ;
        RECT 1093.610 1495.720 1108.410 1496.410 ;
        RECT 1109.250 1495.720 1124.510 1496.410 ;
        RECT 1125.350 1495.720 1140.610 1496.410 ;
        RECT 1141.450 1495.720 1156.250 1496.410 ;
        RECT 1157.090 1495.720 1172.350 1496.410 ;
        RECT 1173.190 1495.720 1188.450 1496.410 ;
        RECT 1189.290 1495.720 1204.090 1496.410 ;
        RECT 1204.930 1495.720 1220.190 1496.410 ;
        RECT 1221.030 1495.720 1236.290 1496.410 ;
        RECT 1237.130 1495.720 1251.930 1496.410 ;
        RECT 1252.770 1495.720 1268.030 1496.410 ;
        RECT 1268.870 1495.720 1284.130 1496.410 ;
        RECT 1284.970 1495.720 1300.230 1496.410 ;
        RECT 1301.070 1495.720 1315.870 1496.410 ;
        RECT 1316.710 1495.720 1331.970 1496.410 ;
        RECT 1332.810 1495.720 1348.070 1496.410 ;
        RECT 1348.910 1495.720 1363.710 1496.410 ;
        RECT 1364.550 1495.720 1379.810 1496.410 ;
        RECT 1380.650 1495.720 1395.910 1496.410 ;
        RECT 1396.750 1495.720 1411.550 1496.410 ;
        RECT 1412.390 1495.720 1427.650 1496.410 ;
        RECT 1428.490 1495.720 1443.750 1496.410 ;
        RECT 1444.590 1495.720 1459.390 1496.410 ;
        RECT 1460.230 1495.720 1475.490 1496.410 ;
        RECT 1476.330 1495.720 1491.590 1496.410 ;
        RECT 6.990 4.280 1492.140 1495.720 ;
        RECT 6.990 3.670 9.010 4.280 ;
        RECT 9.850 3.670 27.410 4.280 ;
        RECT 28.250 3.670 45.810 4.280 ;
        RECT 46.650 3.670 64.210 4.280 ;
        RECT 65.050 3.670 83.070 4.280 ;
        RECT 83.910 3.670 101.470 4.280 ;
        RECT 102.310 3.670 119.870 4.280 ;
        RECT 120.710 3.670 138.270 4.280 ;
        RECT 139.110 3.670 157.130 4.280 ;
        RECT 157.970 3.670 175.530 4.280 ;
        RECT 176.370 3.670 193.930 4.280 ;
        RECT 194.770 3.670 212.330 4.280 ;
        RECT 213.170 3.670 231.190 4.280 ;
        RECT 232.030 3.670 249.590 4.280 ;
        RECT 250.430 3.670 267.990 4.280 ;
        RECT 268.830 3.670 286.390 4.280 ;
        RECT 287.230 3.670 305.250 4.280 ;
        RECT 306.090 3.670 323.650 4.280 ;
        RECT 324.490 3.670 342.050 4.280 ;
        RECT 342.890 3.670 360.450 4.280 ;
        RECT 361.290 3.670 379.310 4.280 ;
        RECT 380.150 3.670 397.710 4.280 ;
        RECT 398.550 3.670 416.110 4.280 ;
        RECT 416.950 3.670 434.510 4.280 ;
        RECT 435.350 3.670 453.370 4.280 ;
        RECT 454.210 3.670 471.770 4.280 ;
        RECT 472.610 3.670 490.170 4.280 ;
        RECT 491.010 3.670 509.030 4.280 ;
        RECT 509.870 3.670 527.430 4.280 ;
        RECT 528.270 3.670 545.830 4.280 ;
        RECT 546.670 3.670 564.230 4.280 ;
        RECT 565.070 3.670 583.090 4.280 ;
        RECT 583.930 3.670 601.490 4.280 ;
        RECT 602.330 3.670 619.890 4.280 ;
        RECT 620.730 3.670 638.290 4.280 ;
        RECT 639.130 3.670 657.150 4.280 ;
        RECT 657.990 3.670 675.550 4.280 ;
        RECT 676.390 3.670 693.950 4.280 ;
        RECT 694.790 3.670 712.350 4.280 ;
        RECT 713.190 3.670 731.210 4.280 ;
        RECT 732.050 3.670 749.610 4.280 ;
        RECT 750.450 3.670 768.010 4.280 ;
        RECT 768.850 3.670 786.410 4.280 ;
        RECT 787.250 3.670 805.270 4.280 ;
        RECT 806.110 3.670 823.670 4.280 ;
        RECT 824.510 3.670 842.070 4.280 ;
        RECT 842.910 3.670 860.470 4.280 ;
        RECT 861.310 3.670 879.330 4.280 ;
        RECT 880.170 3.670 897.730 4.280 ;
        RECT 898.570 3.670 916.130 4.280 ;
        RECT 916.970 3.670 934.530 4.280 ;
        RECT 935.370 3.670 953.390 4.280 ;
        RECT 954.230 3.670 971.790 4.280 ;
        RECT 972.630 3.670 990.190 4.280 ;
        RECT 991.030 3.670 1009.050 4.280 ;
        RECT 1009.890 3.670 1027.450 4.280 ;
        RECT 1028.290 3.670 1045.850 4.280 ;
        RECT 1046.690 3.670 1064.250 4.280 ;
        RECT 1065.090 3.670 1083.110 4.280 ;
        RECT 1083.950 3.670 1101.510 4.280 ;
        RECT 1102.350 3.670 1119.910 4.280 ;
        RECT 1120.750 3.670 1138.310 4.280 ;
        RECT 1139.150 3.670 1157.170 4.280 ;
        RECT 1158.010 3.670 1175.570 4.280 ;
        RECT 1176.410 3.670 1193.970 4.280 ;
        RECT 1194.810 3.670 1212.370 4.280 ;
        RECT 1213.210 3.670 1231.230 4.280 ;
        RECT 1232.070 3.670 1249.630 4.280 ;
        RECT 1250.470 3.670 1268.030 4.280 ;
        RECT 1268.870 3.670 1286.430 4.280 ;
        RECT 1287.270 3.670 1305.290 4.280 ;
        RECT 1306.130 3.670 1323.690 4.280 ;
        RECT 1324.530 3.670 1342.090 4.280 ;
        RECT 1342.930 3.670 1360.490 4.280 ;
        RECT 1361.330 3.670 1379.350 4.280 ;
        RECT 1380.190 3.670 1397.750 4.280 ;
        RECT 1398.590 3.670 1416.150 4.280 ;
        RECT 1416.990 3.670 1434.550 4.280 ;
        RECT 1435.390 3.670 1453.410 4.280 ;
        RECT 1454.250 3.670 1471.810 4.280 ;
        RECT 1472.650 3.670 1490.210 4.280 ;
        RECT 1491.050 3.670 1492.140 4.280 ;
      LAYER met3 ;
        RECT 4.400 1491.600 1496.000 1491.745 ;
        RECT 4.400 1490.880 1495.600 1491.600 ;
        RECT 4.000 1490.200 1495.600 1490.880 ;
        RECT 4.000 1475.960 1496.000 1490.200 ;
        RECT 4.400 1474.560 1496.000 1475.960 ;
        RECT 4.000 1473.240 1496.000 1474.560 ;
        RECT 4.000 1471.840 1495.600 1473.240 ;
        RECT 4.000 1459.640 1496.000 1471.840 ;
        RECT 4.400 1458.240 1496.000 1459.640 ;
        RECT 4.000 1455.560 1496.000 1458.240 ;
        RECT 4.000 1454.160 1495.600 1455.560 ;
        RECT 4.000 1443.320 1496.000 1454.160 ;
        RECT 4.400 1441.920 1496.000 1443.320 ;
        RECT 4.000 1437.200 1496.000 1441.920 ;
        RECT 4.000 1435.800 1495.600 1437.200 ;
        RECT 4.000 1427.000 1496.000 1435.800 ;
        RECT 4.400 1425.600 1496.000 1427.000 ;
        RECT 4.000 1419.520 1496.000 1425.600 ;
        RECT 4.000 1418.120 1495.600 1419.520 ;
        RECT 4.000 1410.680 1496.000 1418.120 ;
        RECT 4.400 1409.280 1496.000 1410.680 ;
        RECT 4.000 1401.160 1496.000 1409.280 ;
        RECT 4.000 1399.760 1495.600 1401.160 ;
        RECT 4.000 1394.360 1496.000 1399.760 ;
        RECT 4.400 1392.960 1496.000 1394.360 ;
        RECT 4.000 1382.800 1496.000 1392.960 ;
        RECT 4.000 1381.400 1495.600 1382.800 ;
        RECT 4.000 1378.040 1496.000 1381.400 ;
        RECT 4.400 1376.640 1496.000 1378.040 ;
        RECT 4.000 1365.120 1496.000 1376.640 ;
        RECT 4.000 1363.720 1495.600 1365.120 ;
        RECT 4.000 1361.720 1496.000 1363.720 ;
        RECT 4.400 1360.320 1496.000 1361.720 ;
        RECT 4.000 1346.760 1496.000 1360.320 ;
        RECT 4.000 1345.400 1495.600 1346.760 ;
        RECT 4.400 1345.360 1495.600 1345.400 ;
        RECT 4.400 1344.000 1496.000 1345.360 ;
        RECT 4.000 1329.080 1496.000 1344.000 ;
        RECT 4.400 1327.680 1495.600 1329.080 ;
        RECT 4.000 1312.760 1496.000 1327.680 ;
        RECT 4.400 1311.360 1496.000 1312.760 ;
        RECT 4.000 1310.720 1496.000 1311.360 ;
        RECT 4.000 1309.320 1495.600 1310.720 ;
        RECT 4.000 1296.440 1496.000 1309.320 ;
        RECT 4.400 1295.040 1496.000 1296.440 ;
        RECT 4.000 1293.040 1496.000 1295.040 ;
        RECT 4.000 1291.640 1495.600 1293.040 ;
        RECT 4.000 1280.120 1496.000 1291.640 ;
        RECT 4.400 1278.720 1496.000 1280.120 ;
        RECT 4.000 1274.680 1496.000 1278.720 ;
        RECT 4.000 1273.280 1495.600 1274.680 ;
        RECT 4.000 1263.800 1496.000 1273.280 ;
        RECT 4.400 1262.400 1496.000 1263.800 ;
        RECT 4.000 1256.320 1496.000 1262.400 ;
        RECT 4.000 1254.920 1495.600 1256.320 ;
        RECT 4.000 1247.480 1496.000 1254.920 ;
        RECT 4.400 1246.080 1496.000 1247.480 ;
        RECT 4.000 1238.640 1496.000 1246.080 ;
        RECT 4.000 1237.240 1495.600 1238.640 ;
        RECT 4.000 1231.160 1496.000 1237.240 ;
        RECT 4.400 1229.760 1496.000 1231.160 ;
        RECT 4.000 1220.280 1496.000 1229.760 ;
        RECT 4.000 1218.880 1495.600 1220.280 ;
        RECT 4.000 1214.840 1496.000 1218.880 ;
        RECT 4.400 1213.440 1496.000 1214.840 ;
        RECT 4.000 1202.600 1496.000 1213.440 ;
        RECT 4.000 1201.200 1495.600 1202.600 ;
        RECT 4.000 1198.520 1496.000 1201.200 ;
        RECT 4.400 1197.120 1496.000 1198.520 ;
        RECT 4.000 1184.240 1496.000 1197.120 ;
        RECT 4.000 1182.840 1495.600 1184.240 ;
        RECT 4.000 1182.200 1496.000 1182.840 ;
        RECT 4.400 1180.800 1496.000 1182.200 ;
        RECT 4.000 1166.560 1496.000 1180.800 ;
        RECT 4.000 1165.880 1495.600 1166.560 ;
        RECT 4.400 1165.160 1495.600 1165.880 ;
        RECT 4.400 1164.480 1496.000 1165.160 ;
        RECT 4.000 1149.560 1496.000 1164.480 ;
        RECT 4.400 1148.200 1496.000 1149.560 ;
        RECT 4.400 1148.160 1495.600 1148.200 ;
        RECT 4.000 1146.800 1495.600 1148.160 ;
        RECT 4.000 1133.240 1496.000 1146.800 ;
        RECT 4.400 1131.840 1496.000 1133.240 ;
        RECT 4.000 1129.840 1496.000 1131.840 ;
        RECT 4.000 1128.440 1495.600 1129.840 ;
        RECT 4.000 1116.920 1496.000 1128.440 ;
        RECT 4.400 1115.520 1496.000 1116.920 ;
        RECT 4.000 1112.160 1496.000 1115.520 ;
        RECT 4.000 1110.760 1495.600 1112.160 ;
        RECT 4.000 1100.600 1496.000 1110.760 ;
        RECT 4.400 1099.200 1496.000 1100.600 ;
        RECT 4.000 1093.800 1496.000 1099.200 ;
        RECT 4.000 1092.400 1495.600 1093.800 ;
        RECT 4.000 1084.280 1496.000 1092.400 ;
        RECT 4.400 1082.880 1496.000 1084.280 ;
        RECT 4.000 1076.120 1496.000 1082.880 ;
        RECT 4.000 1074.720 1495.600 1076.120 ;
        RECT 4.000 1067.960 1496.000 1074.720 ;
        RECT 4.400 1066.560 1496.000 1067.960 ;
        RECT 4.000 1057.760 1496.000 1066.560 ;
        RECT 4.000 1056.360 1495.600 1057.760 ;
        RECT 4.000 1051.640 1496.000 1056.360 ;
        RECT 4.400 1050.240 1496.000 1051.640 ;
        RECT 4.000 1039.400 1496.000 1050.240 ;
        RECT 4.000 1038.000 1495.600 1039.400 ;
        RECT 4.000 1035.320 1496.000 1038.000 ;
        RECT 4.400 1033.920 1496.000 1035.320 ;
        RECT 4.000 1021.720 1496.000 1033.920 ;
        RECT 4.000 1020.320 1495.600 1021.720 ;
        RECT 4.000 1019.000 1496.000 1020.320 ;
        RECT 4.400 1017.600 1496.000 1019.000 ;
        RECT 4.000 1003.360 1496.000 1017.600 ;
        RECT 4.000 1002.680 1495.600 1003.360 ;
        RECT 4.400 1001.960 1495.600 1002.680 ;
        RECT 4.400 1001.280 1496.000 1001.960 ;
        RECT 4.000 986.360 1496.000 1001.280 ;
        RECT 4.400 985.680 1496.000 986.360 ;
        RECT 4.400 984.960 1495.600 985.680 ;
        RECT 4.000 984.280 1495.600 984.960 ;
        RECT 4.000 970.040 1496.000 984.280 ;
        RECT 4.400 968.640 1496.000 970.040 ;
        RECT 4.000 967.320 1496.000 968.640 ;
        RECT 4.000 965.920 1495.600 967.320 ;
        RECT 4.000 953.720 1496.000 965.920 ;
        RECT 4.400 952.320 1496.000 953.720 ;
        RECT 4.000 949.640 1496.000 952.320 ;
        RECT 4.000 948.240 1495.600 949.640 ;
        RECT 4.000 937.400 1496.000 948.240 ;
        RECT 4.400 936.000 1496.000 937.400 ;
        RECT 4.000 931.280 1496.000 936.000 ;
        RECT 4.000 929.880 1495.600 931.280 ;
        RECT 4.000 921.080 1496.000 929.880 ;
        RECT 4.400 919.680 1496.000 921.080 ;
        RECT 4.000 912.920 1496.000 919.680 ;
        RECT 4.000 911.520 1495.600 912.920 ;
        RECT 4.000 904.760 1496.000 911.520 ;
        RECT 4.400 903.360 1496.000 904.760 ;
        RECT 4.000 895.240 1496.000 903.360 ;
        RECT 4.000 893.840 1495.600 895.240 ;
        RECT 4.000 888.440 1496.000 893.840 ;
        RECT 4.400 887.040 1496.000 888.440 ;
        RECT 4.000 876.880 1496.000 887.040 ;
        RECT 4.000 875.480 1495.600 876.880 ;
        RECT 4.000 872.120 1496.000 875.480 ;
        RECT 4.400 870.720 1496.000 872.120 ;
        RECT 4.000 859.200 1496.000 870.720 ;
        RECT 4.000 857.800 1495.600 859.200 ;
        RECT 4.000 855.800 1496.000 857.800 ;
        RECT 4.400 854.400 1496.000 855.800 ;
        RECT 4.000 840.840 1496.000 854.400 ;
        RECT 4.000 839.480 1495.600 840.840 ;
        RECT 4.400 839.440 1495.600 839.480 ;
        RECT 4.400 838.080 1496.000 839.440 ;
        RECT 4.000 823.160 1496.000 838.080 ;
        RECT 4.400 821.760 1495.600 823.160 ;
        RECT 4.000 806.840 1496.000 821.760 ;
        RECT 4.400 805.440 1496.000 806.840 ;
        RECT 4.000 804.800 1496.000 805.440 ;
        RECT 4.000 803.400 1495.600 804.800 ;
        RECT 4.000 790.520 1496.000 803.400 ;
        RECT 4.400 789.120 1496.000 790.520 ;
        RECT 4.000 786.440 1496.000 789.120 ;
        RECT 4.000 785.040 1495.600 786.440 ;
        RECT 4.000 774.200 1496.000 785.040 ;
        RECT 4.400 772.800 1496.000 774.200 ;
        RECT 4.000 768.760 1496.000 772.800 ;
        RECT 4.000 767.360 1495.600 768.760 ;
        RECT 4.000 758.560 1496.000 767.360 ;
        RECT 4.400 757.160 1496.000 758.560 ;
        RECT 4.000 750.400 1496.000 757.160 ;
        RECT 4.000 749.000 1495.600 750.400 ;
        RECT 4.000 742.240 1496.000 749.000 ;
        RECT 4.400 740.840 1496.000 742.240 ;
        RECT 4.000 732.720 1496.000 740.840 ;
        RECT 4.000 731.320 1495.600 732.720 ;
        RECT 4.000 725.920 1496.000 731.320 ;
        RECT 4.400 724.520 1496.000 725.920 ;
        RECT 4.000 714.360 1496.000 724.520 ;
        RECT 4.000 712.960 1495.600 714.360 ;
        RECT 4.000 709.600 1496.000 712.960 ;
        RECT 4.400 708.200 1496.000 709.600 ;
        RECT 4.000 696.000 1496.000 708.200 ;
        RECT 4.000 694.600 1495.600 696.000 ;
        RECT 4.000 693.280 1496.000 694.600 ;
        RECT 4.400 691.880 1496.000 693.280 ;
        RECT 4.000 678.320 1496.000 691.880 ;
        RECT 4.000 676.960 1495.600 678.320 ;
        RECT 4.400 676.920 1495.600 676.960 ;
        RECT 4.400 675.560 1496.000 676.920 ;
        RECT 4.000 660.640 1496.000 675.560 ;
        RECT 4.400 659.960 1496.000 660.640 ;
        RECT 4.400 659.240 1495.600 659.960 ;
        RECT 4.000 658.560 1495.600 659.240 ;
        RECT 4.000 644.320 1496.000 658.560 ;
        RECT 4.400 642.920 1496.000 644.320 ;
        RECT 4.000 642.280 1496.000 642.920 ;
        RECT 4.000 640.880 1495.600 642.280 ;
        RECT 4.000 628.000 1496.000 640.880 ;
        RECT 4.400 626.600 1496.000 628.000 ;
        RECT 4.000 623.920 1496.000 626.600 ;
        RECT 4.000 622.520 1495.600 623.920 ;
        RECT 4.000 611.680 1496.000 622.520 ;
        RECT 4.400 610.280 1496.000 611.680 ;
        RECT 4.000 606.240 1496.000 610.280 ;
        RECT 4.000 604.840 1495.600 606.240 ;
        RECT 4.000 595.360 1496.000 604.840 ;
        RECT 4.400 593.960 1496.000 595.360 ;
        RECT 4.000 587.880 1496.000 593.960 ;
        RECT 4.000 586.480 1495.600 587.880 ;
        RECT 4.000 579.040 1496.000 586.480 ;
        RECT 4.400 577.640 1496.000 579.040 ;
        RECT 4.000 569.520 1496.000 577.640 ;
        RECT 4.000 568.120 1495.600 569.520 ;
        RECT 4.000 562.720 1496.000 568.120 ;
        RECT 4.400 561.320 1496.000 562.720 ;
        RECT 4.000 551.840 1496.000 561.320 ;
        RECT 4.000 550.440 1495.600 551.840 ;
        RECT 4.000 546.400 1496.000 550.440 ;
        RECT 4.400 545.000 1496.000 546.400 ;
        RECT 4.000 533.480 1496.000 545.000 ;
        RECT 4.000 532.080 1495.600 533.480 ;
        RECT 4.000 530.080 1496.000 532.080 ;
        RECT 4.400 528.680 1496.000 530.080 ;
        RECT 4.000 515.800 1496.000 528.680 ;
        RECT 4.000 514.400 1495.600 515.800 ;
        RECT 4.000 513.760 1496.000 514.400 ;
        RECT 4.400 512.360 1496.000 513.760 ;
        RECT 4.000 497.440 1496.000 512.360 ;
        RECT 4.400 496.040 1495.600 497.440 ;
        RECT 4.000 481.120 1496.000 496.040 ;
        RECT 4.400 479.760 1496.000 481.120 ;
        RECT 4.400 479.720 1495.600 479.760 ;
        RECT 4.000 478.360 1495.600 479.720 ;
        RECT 4.000 464.800 1496.000 478.360 ;
        RECT 4.400 463.400 1496.000 464.800 ;
        RECT 4.000 461.400 1496.000 463.400 ;
        RECT 4.000 460.000 1495.600 461.400 ;
        RECT 4.000 448.480 1496.000 460.000 ;
        RECT 4.400 447.080 1496.000 448.480 ;
        RECT 4.000 443.040 1496.000 447.080 ;
        RECT 4.000 441.640 1495.600 443.040 ;
        RECT 4.000 432.160 1496.000 441.640 ;
        RECT 4.400 430.760 1496.000 432.160 ;
        RECT 4.000 425.360 1496.000 430.760 ;
        RECT 4.000 423.960 1495.600 425.360 ;
        RECT 4.000 415.840 1496.000 423.960 ;
        RECT 4.400 414.440 1496.000 415.840 ;
        RECT 4.000 407.000 1496.000 414.440 ;
        RECT 4.000 405.600 1495.600 407.000 ;
        RECT 4.000 399.520 1496.000 405.600 ;
        RECT 4.400 398.120 1496.000 399.520 ;
        RECT 4.000 389.320 1496.000 398.120 ;
        RECT 4.000 387.920 1495.600 389.320 ;
        RECT 4.000 383.200 1496.000 387.920 ;
        RECT 4.400 381.800 1496.000 383.200 ;
        RECT 4.000 370.960 1496.000 381.800 ;
        RECT 4.000 369.560 1495.600 370.960 ;
        RECT 4.000 366.880 1496.000 369.560 ;
        RECT 4.400 365.480 1496.000 366.880 ;
        RECT 4.000 352.600 1496.000 365.480 ;
        RECT 4.000 351.200 1495.600 352.600 ;
        RECT 4.000 350.560 1496.000 351.200 ;
        RECT 4.400 349.160 1496.000 350.560 ;
        RECT 4.000 334.920 1496.000 349.160 ;
        RECT 4.000 334.240 1495.600 334.920 ;
        RECT 4.400 333.520 1495.600 334.240 ;
        RECT 4.400 332.840 1496.000 333.520 ;
        RECT 4.000 317.920 1496.000 332.840 ;
        RECT 4.400 316.560 1496.000 317.920 ;
        RECT 4.400 316.520 1495.600 316.560 ;
        RECT 4.000 315.160 1495.600 316.520 ;
        RECT 4.000 301.600 1496.000 315.160 ;
        RECT 4.400 300.200 1496.000 301.600 ;
        RECT 4.000 298.880 1496.000 300.200 ;
        RECT 4.000 297.480 1495.600 298.880 ;
        RECT 4.000 285.280 1496.000 297.480 ;
        RECT 4.400 283.880 1496.000 285.280 ;
        RECT 4.000 280.520 1496.000 283.880 ;
        RECT 4.000 279.120 1495.600 280.520 ;
        RECT 4.000 268.960 1496.000 279.120 ;
        RECT 4.400 267.560 1496.000 268.960 ;
        RECT 4.000 262.840 1496.000 267.560 ;
        RECT 4.000 261.440 1495.600 262.840 ;
        RECT 4.000 252.640 1496.000 261.440 ;
        RECT 4.400 251.240 1496.000 252.640 ;
        RECT 4.000 244.480 1496.000 251.240 ;
        RECT 4.000 243.080 1495.600 244.480 ;
        RECT 4.000 236.320 1496.000 243.080 ;
        RECT 4.400 234.920 1496.000 236.320 ;
        RECT 4.000 226.120 1496.000 234.920 ;
        RECT 4.000 224.720 1495.600 226.120 ;
        RECT 4.000 220.000 1496.000 224.720 ;
        RECT 4.400 218.600 1496.000 220.000 ;
        RECT 4.000 208.440 1496.000 218.600 ;
        RECT 4.000 207.040 1495.600 208.440 ;
        RECT 4.000 203.680 1496.000 207.040 ;
        RECT 4.400 202.280 1496.000 203.680 ;
        RECT 4.000 190.080 1496.000 202.280 ;
        RECT 4.000 188.680 1495.600 190.080 ;
        RECT 4.000 187.360 1496.000 188.680 ;
        RECT 4.400 185.960 1496.000 187.360 ;
        RECT 4.000 172.400 1496.000 185.960 ;
        RECT 4.000 171.040 1495.600 172.400 ;
        RECT 4.400 171.000 1495.600 171.040 ;
        RECT 4.400 169.640 1496.000 171.000 ;
        RECT 4.000 154.720 1496.000 169.640 ;
        RECT 4.400 154.040 1496.000 154.720 ;
        RECT 4.400 153.320 1495.600 154.040 ;
        RECT 4.000 152.640 1495.600 153.320 ;
        RECT 4.000 138.400 1496.000 152.640 ;
        RECT 4.400 137.000 1496.000 138.400 ;
        RECT 4.000 136.360 1496.000 137.000 ;
        RECT 4.000 134.960 1495.600 136.360 ;
        RECT 4.000 122.080 1496.000 134.960 ;
        RECT 4.400 120.680 1496.000 122.080 ;
        RECT 4.000 118.000 1496.000 120.680 ;
        RECT 4.000 116.600 1495.600 118.000 ;
        RECT 4.000 105.760 1496.000 116.600 ;
        RECT 4.400 104.360 1496.000 105.760 ;
        RECT 4.000 99.640 1496.000 104.360 ;
        RECT 4.000 98.240 1495.600 99.640 ;
        RECT 4.000 89.440 1496.000 98.240 ;
        RECT 4.400 88.040 1496.000 89.440 ;
        RECT 4.000 81.960 1496.000 88.040 ;
        RECT 4.000 80.560 1495.600 81.960 ;
        RECT 4.000 73.120 1496.000 80.560 ;
        RECT 4.400 71.720 1496.000 73.120 ;
        RECT 4.000 63.600 1496.000 71.720 ;
        RECT 4.000 62.200 1495.600 63.600 ;
        RECT 4.000 56.800 1496.000 62.200 ;
        RECT 4.400 55.400 1496.000 56.800 ;
        RECT 4.000 45.920 1496.000 55.400 ;
        RECT 4.000 44.520 1495.600 45.920 ;
        RECT 4.000 40.480 1496.000 44.520 ;
        RECT 4.400 39.080 1496.000 40.480 ;
        RECT 4.000 27.560 1496.000 39.080 ;
        RECT 4.000 26.160 1495.600 27.560 ;
        RECT 4.000 24.160 1496.000 26.160 ;
        RECT 4.400 22.760 1496.000 24.160 ;
        RECT 4.000 9.880 1496.000 22.760 ;
        RECT 4.000 8.520 1495.600 9.880 ;
        RECT 4.400 8.480 1495.600 8.520 ;
        RECT 4.400 7.655 1496.000 8.480 ;
      LAYER met4 ;
        RECT 170.495 11.735 174.240 1486.305 ;
        RECT 176.640 11.735 251.040 1486.305 ;
        RECT 253.440 11.735 327.840 1486.305 ;
        RECT 330.240 11.735 404.640 1486.305 ;
        RECT 407.040 11.735 481.440 1486.305 ;
        RECT 483.840 11.735 558.240 1486.305 ;
        RECT 560.640 11.735 635.040 1486.305 ;
        RECT 637.440 11.735 711.840 1486.305 ;
        RECT 714.240 11.735 788.640 1486.305 ;
        RECT 791.040 11.735 865.440 1486.305 ;
        RECT 867.840 11.735 942.240 1486.305 ;
        RECT 944.640 11.735 989.625 1486.305 ;
  END
END core
END LIBRARY

