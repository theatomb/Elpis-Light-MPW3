VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO regfile
  CLASS BLOCK ;
  FOREIGN regfile ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 450.000 ;
  PIN a[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 102.040 450.000 102.640 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 250.280 450.000 250.880 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 73.480 450.000 74.080 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 446.000 165.050 450.000 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 176.840 450.000 177.440 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 412.120 450.000 412.720 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 446.000 54.650 450.000 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 338.680 450.000 339.280 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 446.000 274.530 450.000 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 446.000 224.850 450.000 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 308.760 450.000 309.360 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 446.000 304.890 450.000 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 446.000 335.250 450.000 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 368.600 450.000 369.200 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 446.000 144.810 450.000 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 446.000 105.250 450.000 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 446.000 325.130 450.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 446.000 4.970 450.000 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END a[9]
  PIN addr_a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END addr_a[0]
  PIN addr_a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 446.000 35.330 450.000 ;
    END
  END addr_a[1]
  PIN addr_a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END addr_a[2]
  PIN addr_a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 280.200 450.000 280.800 ;
    END
  END addr_a[3]
  PIN addr_a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 446.000 444.730 450.000 ;
    END
  END addr_a[4]
  PIN addr_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 28.600 450.000 29.200 ;
    END
  END addr_b[0]
  PIN addr_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END addr_b[1]
  PIN addr_b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END addr_b[2]
  PIN addr_b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 43.560 450.000 44.160 ;
    END
  END addr_b[3]
  PIN addr_b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 117.000 450.000 117.600 ;
    END
  END addr_b[4]
  PIN addr_d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END addr_d[0]
  PIN addr_d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END addr_d[1]
  PIN addr_d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 220.360 450.000 220.960 ;
    END
  END addr_d[2]
  PIN addr_d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 446.000 95.130 450.000 ;
    END
  END addr_d[3]
  PIN addr_d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END addr_d[4]
  PIN b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 446.000 234.970 450.000 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 353.640 450.000 354.240 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 383.560 450.000 384.160 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 446.000 434.610 450.000 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 446.000 195.410 450.000 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 131.960 450.000 132.560 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 446.000 374.810 450.000 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 446.000 315.010 450.000 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 446.000 424.490 450.000 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 446.000 384.930 450.000 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 205.400 450.000 206.000 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 446.000 255.210 450.000 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 446.000 245.090 450.000 ;
    END
  END b[31]
  PIN b[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 446.000 85.010 450.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 442.040 450.000 442.640 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 87.080 450.000 87.680 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END b[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END clk
  PIN d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 293.800 450.000 294.400 ;
    END
  END d[0]
  PIN d[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 446.000 185.290 450.000 ;
    END
  END d[10]
  PIN d[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 446.000 364.690 450.000 ;
    END
  END d[11]
  PIN d[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 446.000 294.770 450.000 ;
    END
  END d[12]
  PIN d[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 446.000 405.170 450.000 ;
    END
  END d[13]
  PIN d[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END d[14]
  PIN d[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END d[15]
  PIN d[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END d[16]
  PIN d[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 446.000 125.490 450.000 ;
    END
  END d[17]
  PIN d[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 446.000 214.730 450.000 ;
    END
  END d[18]
  PIN d[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 146.920 450.000 147.520 ;
    END
  END d[19]
  PIN d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 446.000 204.610 450.000 ;
    END
  END d[1]
  PIN d[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END d[20]
  PIN d[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 446.000 115.370 450.000 ;
    END
  END d[21]
  PIN d[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END d[22]
  PIN d[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END d[23]
  PIN d[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 446.000 64.770 450.000 ;
    END
  END d[24]
  PIN d[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END d[25]
  PIN d[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END d[26]
  PIN d[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 446.000 45.450 450.000 ;
    END
  END d[27]
  PIN d[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 446.000 414.370 450.000 ;
    END
  END d[28]
  PIN d[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END d[29]
  PIN d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 13.640 450.000 14.240 ;
    END
  END d[2]
  PIN d[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END d[30]
  PIN d[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END d[31]
  PIN d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 446.000 175.170 450.000 ;
    END
  END d[3]
  PIN d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END d[4]
  PIN d[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END d[5]
  PIN d[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END d[6]
  PIN d[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END d[7]
  PIN d[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 323.720 450.000 324.320 ;
    END
  END d[8]
  PIN d[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 190.440 450.000 191.040 ;
    END
  END d[9]
  PIN dest_read[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END dest_read[0]
  PIN dest_read[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END dest_read[1]
  PIN dest_read[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 58.520 450.000 59.120 ;
    END
  END dest_read[2]
  PIN dest_read[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END dest_read[3]
  PIN dest_read[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 235.320 450.000 235.920 ;
    END
  END dest_read[4]
  PIN dest_value[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 397.160 450.000 397.760 ;
    END
  END dest_value[0]
  PIN dest_value[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END dest_value[10]
  PIN dest_value[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 427.080 450.000 427.680 ;
    END
  END dest_value[11]
  PIN dest_value[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END dest_value[12]
  PIN dest_value[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END dest_value[13]
  PIN dest_value[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END dest_value[14]
  PIN dest_value[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END dest_value[15]
  PIN dest_value[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END dest_value[16]
  PIN dest_value[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END dest_value[17]
  PIN dest_value[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 446.000 154.930 450.000 ;
    END
  END dest_value[18]
  PIN dest_value[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 446.000 284.650 450.000 ;
    END
  END dest_value[19]
  PIN dest_value[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END dest_value[1]
  PIN dest_value[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END dest_value[20]
  PIN dest_value[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END dest_value[21]
  PIN dest_value[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END dest_value[22]
  PIN dest_value[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 446.000 265.330 450.000 ;
    END
  END dest_value[23]
  PIN dest_value[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END dest_value[24]
  PIN dest_value[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 446.000 395.050 450.000 ;
    END
  END dest_value[25]
  PIN dest_value[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END dest_value[26]
  PIN dest_value[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 446.000 25.210 450.000 ;
    END
  END dest_value[27]
  PIN dest_value[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END dest_value[28]
  PIN dest_value[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END dest_value[29]
  PIN dest_value[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END dest_value[2]
  PIN dest_value[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END dest_value[30]
  PIN dest_value[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 265.240 450.000 265.840 ;
    END
  END dest_value[31]
  PIN dest_value[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END dest_value[3]
  PIN dest_value[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 446.000 354.570 450.000 ;
    END
  END dest_value[4]
  PIN dest_value[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 446.000 344.450 450.000 ;
    END
  END dest_value[5]
  PIN dest_value[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 446.000 74.890 450.000 ;
    END
  END dest_value[6]
  PIN dest_value[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 446.000 134.690 450.000 ;
    END
  END dest_value[7]
  PIN dest_value[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END dest_value[8]
  PIN dest_value[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END dest_value[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 446.000 15.090 450.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 438.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 438.160 ;
    END
  END vssd1
  PIN wrd
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 161.880 450.000 162.480 ;
    END
  END wrd
  OBS
      LAYER li1 ;
        RECT 5.520 7.905 444.360 438.005 ;
      LAYER met1 ;
        RECT 0.070 7.520 449.350 438.900 ;
      LAYER met2 ;
        RECT 0.100 445.720 4.410 446.490 ;
        RECT 5.250 445.720 14.530 446.490 ;
        RECT 15.370 445.720 24.650 446.490 ;
        RECT 25.490 445.720 34.770 446.490 ;
        RECT 35.610 445.720 44.890 446.490 ;
        RECT 45.730 445.720 54.090 446.490 ;
        RECT 54.930 445.720 64.210 446.490 ;
        RECT 65.050 445.720 74.330 446.490 ;
        RECT 75.170 445.720 84.450 446.490 ;
        RECT 85.290 445.720 94.570 446.490 ;
        RECT 95.410 445.720 104.690 446.490 ;
        RECT 105.530 445.720 114.810 446.490 ;
        RECT 115.650 445.720 124.930 446.490 ;
        RECT 125.770 445.720 134.130 446.490 ;
        RECT 134.970 445.720 144.250 446.490 ;
        RECT 145.090 445.720 154.370 446.490 ;
        RECT 155.210 445.720 164.490 446.490 ;
        RECT 165.330 445.720 174.610 446.490 ;
        RECT 175.450 445.720 184.730 446.490 ;
        RECT 185.570 445.720 194.850 446.490 ;
        RECT 195.690 445.720 204.050 446.490 ;
        RECT 204.890 445.720 214.170 446.490 ;
        RECT 215.010 445.720 224.290 446.490 ;
        RECT 225.130 445.720 234.410 446.490 ;
        RECT 235.250 445.720 244.530 446.490 ;
        RECT 245.370 445.720 254.650 446.490 ;
        RECT 255.490 445.720 264.770 446.490 ;
        RECT 265.610 445.720 273.970 446.490 ;
        RECT 274.810 445.720 284.090 446.490 ;
        RECT 284.930 445.720 294.210 446.490 ;
        RECT 295.050 445.720 304.330 446.490 ;
        RECT 305.170 445.720 314.450 446.490 ;
        RECT 315.290 445.720 324.570 446.490 ;
        RECT 325.410 445.720 334.690 446.490 ;
        RECT 335.530 445.720 343.890 446.490 ;
        RECT 344.730 445.720 354.010 446.490 ;
        RECT 354.850 445.720 364.130 446.490 ;
        RECT 364.970 445.720 374.250 446.490 ;
        RECT 375.090 445.720 384.370 446.490 ;
        RECT 385.210 445.720 394.490 446.490 ;
        RECT 395.330 445.720 404.610 446.490 ;
        RECT 405.450 445.720 413.810 446.490 ;
        RECT 414.650 445.720 423.930 446.490 ;
        RECT 424.770 445.720 434.050 446.490 ;
        RECT 434.890 445.720 444.170 446.490 ;
        RECT 445.010 445.720 449.320 446.490 ;
        RECT 0.100 4.280 449.320 445.720 ;
        RECT 0.650 3.670 9.010 4.280 ;
        RECT 9.850 3.670 19.130 4.280 ;
        RECT 19.970 3.670 29.250 4.280 ;
        RECT 30.090 3.670 39.370 4.280 ;
        RECT 40.210 3.670 49.490 4.280 ;
        RECT 50.330 3.670 59.610 4.280 ;
        RECT 60.450 3.670 69.730 4.280 ;
        RECT 70.570 3.670 78.930 4.280 ;
        RECT 79.770 3.670 89.050 4.280 ;
        RECT 89.890 3.670 99.170 4.280 ;
        RECT 100.010 3.670 109.290 4.280 ;
        RECT 110.130 3.670 119.410 4.280 ;
        RECT 120.250 3.670 129.530 4.280 ;
        RECT 130.370 3.670 139.650 4.280 ;
        RECT 140.490 3.670 148.850 4.280 ;
        RECT 149.690 3.670 158.970 4.280 ;
        RECT 159.810 3.670 169.090 4.280 ;
        RECT 169.930 3.670 179.210 4.280 ;
        RECT 180.050 3.670 189.330 4.280 ;
        RECT 190.170 3.670 199.450 4.280 ;
        RECT 200.290 3.670 209.570 4.280 ;
        RECT 210.410 3.670 218.770 4.280 ;
        RECT 219.610 3.670 228.890 4.280 ;
        RECT 229.730 3.670 239.010 4.280 ;
        RECT 239.850 3.670 249.130 4.280 ;
        RECT 249.970 3.670 259.250 4.280 ;
        RECT 260.090 3.670 269.370 4.280 ;
        RECT 270.210 3.670 279.490 4.280 ;
        RECT 280.330 3.670 288.690 4.280 ;
        RECT 289.530 3.670 298.810 4.280 ;
        RECT 299.650 3.670 308.930 4.280 ;
        RECT 309.770 3.670 319.050 4.280 ;
        RECT 319.890 3.670 329.170 4.280 ;
        RECT 330.010 3.670 339.290 4.280 ;
        RECT 340.130 3.670 349.410 4.280 ;
        RECT 350.250 3.670 358.610 4.280 ;
        RECT 359.450 3.670 368.730 4.280 ;
        RECT 369.570 3.670 378.850 4.280 ;
        RECT 379.690 3.670 388.970 4.280 ;
        RECT 389.810 3.670 399.090 4.280 ;
        RECT 399.930 3.670 409.210 4.280 ;
        RECT 410.050 3.670 419.330 4.280 ;
        RECT 420.170 3.670 429.450 4.280 ;
        RECT 430.290 3.670 438.650 4.280 ;
        RECT 439.490 3.670 448.770 4.280 ;
      LAYER met3 ;
        RECT 4.400 441.640 445.600 442.505 ;
        RECT 4.000 428.080 446.000 441.640 ;
        RECT 4.400 426.680 445.600 428.080 ;
        RECT 4.000 414.480 446.000 426.680 ;
        RECT 4.400 413.120 446.000 414.480 ;
        RECT 4.400 413.080 445.600 413.120 ;
        RECT 4.000 411.720 445.600 413.080 ;
        RECT 4.000 399.520 446.000 411.720 ;
        RECT 4.400 398.160 446.000 399.520 ;
        RECT 4.400 398.120 445.600 398.160 ;
        RECT 4.000 396.760 445.600 398.120 ;
        RECT 4.000 384.560 446.000 396.760 ;
        RECT 4.400 383.160 445.600 384.560 ;
        RECT 4.000 369.600 446.000 383.160 ;
        RECT 4.400 368.200 445.600 369.600 ;
        RECT 4.000 354.640 446.000 368.200 ;
        RECT 4.400 353.240 445.600 354.640 ;
        RECT 4.000 339.680 446.000 353.240 ;
        RECT 4.400 338.280 445.600 339.680 ;
        RECT 4.000 324.720 446.000 338.280 ;
        RECT 4.400 323.320 445.600 324.720 ;
        RECT 4.000 311.120 446.000 323.320 ;
        RECT 4.400 309.760 446.000 311.120 ;
        RECT 4.400 309.720 445.600 309.760 ;
        RECT 4.000 308.360 445.600 309.720 ;
        RECT 4.000 296.160 446.000 308.360 ;
        RECT 4.400 294.800 446.000 296.160 ;
        RECT 4.400 294.760 445.600 294.800 ;
        RECT 4.000 293.400 445.600 294.760 ;
        RECT 4.000 281.200 446.000 293.400 ;
        RECT 4.400 279.800 445.600 281.200 ;
        RECT 4.000 266.240 446.000 279.800 ;
        RECT 4.400 264.840 445.600 266.240 ;
        RECT 4.000 251.280 446.000 264.840 ;
        RECT 4.400 249.880 445.600 251.280 ;
        RECT 4.000 236.320 446.000 249.880 ;
        RECT 4.400 234.920 445.600 236.320 ;
        RECT 4.000 221.360 446.000 234.920 ;
        RECT 4.400 219.960 445.600 221.360 ;
        RECT 4.000 207.760 446.000 219.960 ;
        RECT 4.400 206.400 446.000 207.760 ;
        RECT 4.400 206.360 445.600 206.400 ;
        RECT 4.000 205.000 445.600 206.360 ;
        RECT 4.000 192.800 446.000 205.000 ;
        RECT 4.400 191.440 446.000 192.800 ;
        RECT 4.400 191.400 445.600 191.440 ;
        RECT 4.000 190.040 445.600 191.400 ;
        RECT 4.000 177.840 446.000 190.040 ;
        RECT 4.400 176.440 445.600 177.840 ;
        RECT 4.000 162.880 446.000 176.440 ;
        RECT 4.400 161.480 445.600 162.880 ;
        RECT 4.000 147.920 446.000 161.480 ;
        RECT 4.400 146.520 445.600 147.920 ;
        RECT 4.000 132.960 446.000 146.520 ;
        RECT 4.400 131.560 445.600 132.960 ;
        RECT 4.000 118.000 446.000 131.560 ;
        RECT 4.400 116.600 445.600 118.000 ;
        RECT 4.000 104.400 446.000 116.600 ;
        RECT 4.400 103.040 446.000 104.400 ;
        RECT 4.400 103.000 445.600 103.040 ;
        RECT 4.000 101.640 445.600 103.000 ;
        RECT 4.000 89.440 446.000 101.640 ;
        RECT 4.400 88.080 446.000 89.440 ;
        RECT 4.400 88.040 445.600 88.080 ;
        RECT 4.000 86.680 445.600 88.040 ;
        RECT 4.000 74.480 446.000 86.680 ;
        RECT 4.400 73.080 445.600 74.480 ;
        RECT 4.000 59.520 446.000 73.080 ;
        RECT 4.400 58.120 445.600 59.520 ;
        RECT 4.000 44.560 446.000 58.120 ;
        RECT 4.400 43.160 445.600 44.560 ;
        RECT 4.000 29.600 446.000 43.160 ;
        RECT 4.400 28.200 445.600 29.600 ;
        RECT 4.000 14.640 446.000 28.200 ;
        RECT 4.400 13.240 445.600 14.640 ;
        RECT 4.000 10.715 446.000 13.240 ;
      LAYER met4 ;
        RECT 46.295 11.735 97.440 435.705 ;
        RECT 99.840 11.735 174.240 435.705 ;
        RECT 176.640 11.735 251.040 435.705 ;
        RECT 253.440 11.735 327.840 435.705 ;
        RECT 330.240 11.735 404.640 435.705 ;
        RECT 407.040 11.735 440.385 435.705 ;
  END
END regfile
END LIBRARY

