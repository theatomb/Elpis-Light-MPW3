VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO io_output_arbiter
  CLASS BLOCK ;
  FOREIGN io_output_arbiter ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 75.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END clk
  PIN data_core0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END data_core0[0]
  PIN data_core0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 28.600 75.000 29.200 ;
    END
  END data_core0[10]
  PIN data_core0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 71.000 17.850 75.000 ;
    END
  END data_core0[11]
  PIN data_core0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 71.000 21.530 75.000 ;
    END
  END data_core0[12]
  PIN data_core0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END data_core0[13]
  PIN data_core0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 71.000 25.670 75.000 ;
    END
  END data_core0[14]
  PIN data_core0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 71.000 29.810 75.000 ;
    END
  END data_core0[15]
  PIN data_core0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 35.400 75.000 36.000 ;
    END
  END data_core0[16]
  PIN data_core0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END data_core0[17]
  PIN data_core0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END data_core0[18]
  PIN data_core0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 45.600 75.000 46.200 ;
    END
  END data_core0[19]
  PIN data_core0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 4.800 75.000 5.400 ;
    END
  END data_core0[1]
  PIN data_core0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END data_core0[20]
  PIN data_core0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END data_core0[21]
  PIN data_core0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 71.000 41.310 75.000 ;
    END
  END data_core0[22]
  PIN data_core0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 55.800 75.000 56.400 ;
    END
  END data_core0[23]
  PIN data_core0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 71.000 45.450 75.000 ;
    END
  END data_core0[24]
  PIN data_core0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 71.000 53.270 75.000 ;
    END
  END data_core0[25]
  PIN data_core0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END data_core0[26]
  PIN data_core0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 66.000 75.000 66.600 ;
    END
  END data_core0[27]
  PIN data_core0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END data_core0[28]
  PIN data_core0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 71.000 61.090 75.000 ;
    END
  END data_core0[29]
  PIN data_core0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END data_core0[2]
  PIN data_core0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 71.000 65.230 75.000 ;
    END
  END data_core0[30]
  PIN data_core0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 71.000 73.050 75.000 ;
    END
  END data_core0[31]
  PIN data_core0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END data_core0[3]
  PIN data_core0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 11.600 75.000 12.200 ;
    END
  END data_core0[4]
  PIN data_core0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 15.000 75.000 15.600 ;
    END
  END data_core0[5]
  PIN data_core0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END data_core0[6]
  PIN data_core0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 71.000 10.030 75.000 ;
    END
  END data_core0[7]
  PIN data_core0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END data_core0[8]
  PIN data_core0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 71.000 13.710 75.000 ;
    END
  END data_core0[9]
  PIN is_ready_core0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END is_ready_core0
  PIN print_hex_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END print_hex_enable
  PIN print_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 1.400 75.000 2.000 ;
    END
  END print_output[0]
  PIN print_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END print_output[10]
  PIN print_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END print_output[11]
  PIN print_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 32.000 75.000 32.600 ;
    END
  END print_output[12]
  PIN print_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END print_output[13]
  PIN print_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END print_output[14]
  PIN print_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 71.000 33.490 75.000 ;
    END
  END print_output[15]
  PIN print_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 38.800 75.000 39.400 ;
    END
  END print_output[16]
  PIN print_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 71.000 37.630 75.000 ;
    END
  END print_output[17]
  PIN print_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 42.200 75.000 42.800 ;
    END
  END print_output[18]
  PIN print_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END print_output[19]
  PIN print_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 8.200 75.000 8.800 ;
    END
  END print_output[1]
  PIN print_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 49.000 75.000 49.600 ;
    END
  END print_output[20]
  PIN print_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 52.400 75.000 53.000 ;
    END
  END print_output[21]
  PIN print_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END print_output[22]
  PIN print_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END print_output[23]
  PIN print_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 71.000 49.130 75.000 ;
    END
  END print_output[24]
  PIN print_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 59.200 75.000 59.800 ;
    END
  END print_output[25]
  PIN print_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 62.600 75.000 63.200 ;
    END
  END print_output[26]
  PIN print_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 69.400 75.000 70.000 ;
    END
  END print_output[27]
  PIN print_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 71.000 57.410 75.000 ;
    END
  END print_output[28]
  PIN print_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END print_output[29]
  PIN print_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END print_output[2]
  PIN print_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 71.000 68.910 75.000 ;
    END
  END print_output[30]
  PIN print_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 72.800 75.000 73.400 ;
    END
  END print_output[31]
  PIN print_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 71.000 2.210 75.000 ;
    END
  END print_output[3]
  PIN print_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 71.000 5.890 75.000 ;
    END
  END print_output[4]
  PIN print_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 18.400 75.000 19.000 ;
    END
  END print_output[5]
  PIN print_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 21.800 75.000 22.400 ;
    END
  END print_output[6]
  PIN print_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END print_output[7]
  PIN print_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 25.200 75.000 25.800 ;
    END
  END print_output[8]
  PIN print_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END print_output[9]
  PIN req_core0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END req_core0
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.380 10.640 16.980 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.700 10.640 38.300 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.020 10.640 59.620 62.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.040 10.640 27.640 62.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.360 10.640 48.960 62.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 1.785 70.235 62.645 ;
      LAYER met1 ;
        RECT 1.910 1.740 73.070 62.800 ;
      LAYER met2 ;
        RECT 2.490 70.720 5.330 73.285 ;
        RECT 6.170 70.720 9.470 73.285 ;
        RECT 10.310 70.720 13.150 73.285 ;
        RECT 13.990 70.720 17.290 73.285 ;
        RECT 18.130 70.720 20.970 73.285 ;
        RECT 21.810 70.720 25.110 73.285 ;
        RECT 25.950 70.720 29.250 73.285 ;
        RECT 30.090 70.720 32.930 73.285 ;
        RECT 33.770 70.720 37.070 73.285 ;
        RECT 37.910 70.720 40.750 73.285 ;
        RECT 41.590 70.720 44.890 73.285 ;
        RECT 45.730 70.720 48.570 73.285 ;
        RECT 49.410 70.720 52.710 73.285 ;
        RECT 53.550 70.720 56.850 73.285 ;
        RECT 57.690 70.720 60.530 73.285 ;
        RECT 61.370 70.720 64.670 73.285 ;
        RECT 65.510 70.720 68.350 73.285 ;
        RECT 69.190 70.720 72.490 73.285 ;
        RECT 1.940 4.280 73.040 70.720 ;
        RECT 1.940 1.515 2.110 4.280 ;
        RECT 2.950 1.515 6.710 4.280 ;
        RECT 7.550 1.515 11.310 4.280 ;
        RECT 12.150 1.515 15.910 4.280 ;
        RECT 16.750 1.515 20.510 4.280 ;
        RECT 21.350 1.515 25.110 4.280 ;
        RECT 25.950 1.515 30.170 4.280 ;
        RECT 31.010 1.515 34.770 4.280 ;
        RECT 35.610 1.515 39.370 4.280 ;
        RECT 40.210 1.515 43.970 4.280 ;
        RECT 44.810 1.515 48.570 4.280 ;
        RECT 49.410 1.515 53.630 4.280 ;
        RECT 54.470 1.515 58.230 4.280 ;
        RECT 59.070 1.515 62.830 4.280 ;
        RECT 63.670 1.515 67.430 4.280 ;
        RECT 68.270 1.515 72.030 4.280 ;
        RECT 72.870 1.515 73.040 4.280 ;
      LAYER met3 ;
        RECT 4.000 72.400 70.600 73.265 ;
        RECT 4.000 71.760 71.000 72.400 ;
        RECT 4.400 70.400 71.000 71.760 ;
        RECT 4.400 70.360 70.600 70.400 ;
        RECT 4.000 69.000 70.600 70.360 ;
        RECT 4.000 67.000 71.000 69.000 ;
        RECT 4.000 65.640 70.600 67.000 ;
        RECT 4.400 65.600 70.600 65.640 ;
        RECT 4.400 64.240 71.000 65.600 ;
        RECT 4.000 63.600 71.000 64.240 ;
        RECT 4.000 62.200 70.600 63.600 ;
        RECT 4.000 60.200 71.000 62.200 ;
        RECT 4.000 59.520 70.600 60.200 ;
        RECT 4.400 58.800 70.600 59.520 ;
        RECT 4.400 58.120 71.000 58.800 ;
        RECT 4.000 56.800 71.000 58.120 ;
        RECT 4.000 55.400 70.600 56.800 ;
        RECT 4.000 53.400 71.000 55.400 ;
        RECT 4.400 52.000 70.600 53.400 ;
        RECT 4.000 50.000 71.000 52.000 ;
        RECT 4.000 48.600 70.600 50.000 ;
        RECT 4.000 47.280 71.000 48.600 ;
        RECT 4.400 46.600 71.000 47.280 ;
        RECT 4.400 45.880 70.600 46.600 ;
        RECT 4.000 45.200 70.600 45.880 ;
        RECT 4.000 43.200 71.000 45.200 ;
        RECT 4.000 41.800 70.600 43.200 ;
        RECT 4.000 41.160 71.000 41.800 ;
        RECT 4.400 39.800 71.000 41.160 ;
        RECT 4.400 39.760 70.600 39.800 ;
        RECT 4.000 38.400 70.600 39.760 ;
        RECT 4.000 36.400 71.000 38.400 ;
        RECT 4.000 35.000 70.600 36.400 ;
        RECT 4.000 34.360 71.000 35.000 ;
        RECT 4.400 33.000 71.000 34.360 ;
        RECT 4.400 32.960 70.600 33.000 ;
        RECT 4.000 31.600 70.600 32.960 ;
        RECT 4.000 29.600 71.000 31.600 ;
        RECT 4.000 28.240 70.600 29.600 ;
        RECT 4.400 28.200 70.600 28.240 ;
        RECT 4.400 26.840 71.000 28.200 ;
        RECT 4.000 26.200 71.000 26.840 ;
        RECT 4.000 24.800 70.600 26.200 ;
        RECT 4.000 22.800 71.000 24.800 ;
        RECT 4.000 22.120 70.600 22.800 ;
        RECT 4.400 21.400 70.600 22.120 ;
        RECT 4.400 20.720 71.000 21.400 ;
        RECT 4.000 19.400 71.000 20.720 ;
        RECT 4.000 18.000 70.600 19.400 ;
        RECT 4.000 16.000 71.000 18.000 ;
        RECT 4.400 14.600 70.600 16.000 ;
        RECT 4.000 12.600 71.000 14.600 ;
        RECT 4.000 11.200 70.600 12.600 ;
        RECT 4.000 9.880 71.000 11.200 ;
        RECT 4.400 9.200 71.000 9.880 ;
        RECT 4.400 8.480 70.600 9.200 ;
        RECT 4.000 7.800 70.600 8.480 ;
        RECT 4.000 5.800 71.000 7.800 ;
        RECT 4.000 4.400 70.600 5.800 ;
        RECT 4.000 3.760 71.000 4.400 ;
        RECT 4.400 2.400 71.000 3.760 ;
        RECT 4.400 2.360 70.600 2.400 ;
        RECT 4.000 1.535 70.600 2.360 ;
  END
END io_output_arbiter
END LIBRARY

