* NGSPICE file created from sram_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

.subckt sram_wrapper addr0_to_sram[0] addr0_to_sram[10] addr0_to_sram[11] addr0_to_sram[12]
+ addr0_to_sram[13] addr0_to_sram[14] addr0_to_sram[15] addr0_to_sram[16] addr0_to_sram[17]
+ addr0_to_sram[18] addr0_to_sram[19] addr0_to_sram[1] addr0_to_sram[2] addr0_to_sram[3]
+ addr0_to_sram[4] addr0_to_sram[5] addr0_to_sram[6] addr0_to_sram[7] addr0_to_sram[8]
+ addr0_to_sram[9] addr_in[0] addr_in[10] addr_in[11] addr_in[12] addr_in[13] addr_in[14]
+ addr_in[15] addr_in[16] addr_in[17] addr_in[18] addr_in[19] addr_in[1] addr_in[2]
+ addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in[8] addr_in[9] addr_to_core_mem[0]
+ addr_to_core_mem[10] addr_to_core_mem[11] addr_to_core_mem[12] addr_to_core_mem[13]
+ addr_to_core_mem[14] addr_to_core_mem[15] addr_to_core_mem[16] addr_to_core_mem[17]
+ addr_to_core_mem[18] addr_to_core_mem[19] addr_to_core_mem[1] addr_to_core_mem[2]
+ addr_to_core_mem[3] addr_to_core_mem[4] addr_to_core_mem[5] addr_to_core_mem[6]
+ addr_to_core_mem[7] addr_to_core_mem[8] addr_to_core_mem[9] clk csb0_to_sram data_to_core_mem[0]
+ data_to_core_mem[10] data_to_core_mem[11] data_to_core_mem[12] data_to_core_mem[13]
+ data_to_core_mem[14] data_to_core_mem[15] data_to_core_mem[16] data_to_core_mem[17]
+ data_to_core_mem[18] data_to_core_mem[19] data_to_core_mem[1] data_to_core_mem[20]
+ data_to_core_mem[21] data_to_core_mem[22] data_to_core_mem[23] data_to_core_mem[24]
+ data_to_core_mem[25] data_to_core_mem[26] data_to_core_mem[27] data_to_core_mem[28]
+ data_to_core_mem[29] data_to_core_mem[2] data_to_core_mem[30] data_to_core_mem[31]
+ data_to_core_mem[3] data_to_core_mem[4] data_to_core_mem[5] data_to_core_mem[6]
+ data_to_core_mem[7] data_to_core_mem[8] data_to_core_mem[9] din0_to_sram[0] din0_to_sram[10]
+ din0_to_sram[11] din0_to_sram[12] din0_to_sram[13] din0_to_sram[14] din0_to_sram[15]
+ din0_to_sram[16] din0_to_sram[17] din0_to_sram[18] din0_to_sram[19] din0_to_sram[1]
+ din0_to_sram[20] din0_to_sram[21] din0_to_sram[22] din0_to_sram[23] din0_to_sram[24]
+ din0_to_sram[25] din0_to_sram[26] din0_to_sram[27] din0_to_sram[28] din0_to_sram[29]
+ din0_to_sram[2] din0_to_sram[30] din0_to_sram[31] din0_to_sram[3] din0_to_sram[4]
+ din0_to_sram[5] din0_to_sram[6] din0_to_sram[7] din0_to_sram[8] din0_to_sram[9]
+ dout0_to_sram[0] dout0_to_sram[10] dout0_to_sram[11] dout0_to_sram[12] dout0_to_sram[13]
+ dout0_to_sram[14] dout0_to_sram[15] dout0_to_sram[16] dout0_to_sram[17] dout0_to_sram[18]
+ dout0_to_sram[19] dout0_to_sram[1] dout0_to_sram[20] dout0_to_sram[21] dout0_to_sram[22]
+ dout0_to_sram[23] dout0_to_sram[24] dout0_to_sram[25] dout0_to_sram[26] dout0_to_sram[27]
+ dout0_to_sram[28] dout0_to_sram[29] dout0_to_sram[2] dout0_to_sram[30] dout0_to_sram[31]
+ dout0_to_sram[3] dout0_to_sram[4] dout0_to_sram[5] dout0_to_sram[6] dout0_to_sram[7]
+ dout0_to_sram[8] dout0_to_sram[9] is_loading_memory_into_core rd_data_out[0] rd_data_out[100]
+ rd_data_out[101] rd_data_out[102] rd_data_out[103] rd_data_out[104] rd_data_out[105]
+ rd_data_out[106] rd_data_out[107] rd_data_out[108] rd_data_out[109] rd_data_out[10]
+ rd_data_out[110] rd_data_out[111] rd_data_out[112] rd_data_out[113] rd_data_out[114]
+ rd_data_out[115] rd_data_out[116] rd_data_out[117] rd_data_out[118] rd_data_out[119]
+ rd_data_out[11] rd_data_out[120] rd_data_out[121] rd_data_out[122] rd_data_out[123]
+ rd_data_out[124] rd_data_out[125] rd_data_out[126] rd_data_out[127] rd_data_out[12]
+ rd_data_out[13] rd_data_out[14] rd_data_out[15] rd_data_out[16] rd_data_out[17]
+ rd_data_out[18] rd_data_out[19] rd_data_out[1] rd_data_out[20] rd_data_out[21] rd_data_out[22]
+ rd_data_out[23] rd_data_out[24] rd_data_out[25] rd_data_out[26] rd_data_out[27]
+ rd_data_out[28] rd_data_out[29] rd_data_out[2] rd_data_out[30] rd_data_out[31] rd_data_out[32]
+ rd_data_out[33] rd_data_out[34] rd_data_out[35] rd_data_out[36] rd_data_out[37]
+ rd_data_out[38] rd_data_out[39] rd_data_out[3] rd_data_out[40] rd_data_out[41] rd_data_out[42]
+ rd_data_out[43] rd_data_out[44] rd_data_out[45] rd_data_out[46] rd_data_out[47]
+ rd_data_out[48] rd_data_out[49] rd_data_out[4] rd_data_out[50] rd_data_out[51] rd_data_out[52]
+ rd_data_out[53] rd_data_out[54] rd_data_out[55] rd_data_out[56] rd_data_out[57]
+ rd_data_out[58] rd_data_out[59] rd_data_out[5] rd_data_out[60] rd_data_out[61] rd_data_out[62]
+ rd_data_out[63] rd_data_out[64] rd_data_out[65] rd_data_out[66] rd_data_out[67]
+ rd_data_out[68] rd_data_out[69] rd_data_out[6] rd_data_out[70] rd_data_out[71] rd_data_out[72]
+ rd_data_out[73] rd_data_out[74] rd_data_out[75] rd_data_out[76] rd_data_out[77]
+ rd_data_out[78] rd_data_out[79] rd_data_out[7] rd_data_out[80] rd_data_out[81] rd_data_out[82]
+ rd_data_out[83] rd_data_out[84] rd_data_out[85] rd_data_out[86] rd_data_out[87]
+ rd_data_out[88] rd_data_out[89] rd_data_out[8] rd_data_out[90] rd_data_out[91] rd_data_out[92]
+ rd_data_out[93] rd_data_out[94] rd_data_out[95] rd_data_out[96] rd_data_out[97]
+ rd_data_out[98] rd_data_out[99] rd_data_out[9] ready requested reset reset_mem_req
+ spare_wen0_to_sram vccd1 vssd1 we we_to_sram wr_data[0] wr_data[100] wr_data[101]
+ wr_data[102] wr_data[103] wr_data[104] wr_data[105] wr_data[106] wr_data[107] wr_data[108]
+ wr_data[109] wr_data[10] wr_data[110] wr_data[111] wr_data[112] wr_data[113] wr_data[114]
+ wr_data[115] wr_data[116] wr_data[117] wr_data[118] wr_data[119] wr_data[11] wr_data[120]
+ wr_data[121] wr_data[122] wr_data[123] wr_data[124] wr_data[125] wr_data[126] wr_data[127]
+ wr_data[12] wr_data[13] wr_data[14] wr_data[15] wr_data[16] wr_data[17] wr_data[18]
+ wr_data[19] wr_data[1] wr_data[20] wr_data[21] wr_data[22] wr_data[23] wr_data[24]
+ wr_data[25] wr_data[26] wr_data[27] wr_data[28] wr_data[29] wr_data[2] wr_data[30]
+ wr_data[31] wr_data[32] wr_data[33] wr_data[34] wr_data[35] wr_data[36] wr_data[37]
+ wr_data[38] wr_data[39] wr_data[3] wr_data[40] wr_data[41] wr_data[42] wr_data[43]
+ wr_data[44] wr_data[45] wr_data[46] wr_data[47] wr_data[48] wr_data[49] wr_data[4]
+ wr_data[50] wr_data[51] wr_data[52] wr_data[53] wr_data[54] wr_data[55] wr_data[56]
+ wr_data[57] wr_data[58] wr_data[59] wr_data[5] wr_data[60] wr_data[61] wr_data[62]
+ wr_data[63] wr_data[64] wr_data[65] wr_data[66] wr_data[67] wr_data[68] wr_data[69]
+ wr_data[6] wr_data[70] wr_data[71] wr_data[72] wr_data[73] wr_data[74] wr_data[75]
+ wr_data[76] wr_data[77] wr_data[78] wr_data[79] wr_data[7] wr_data[80] wr_data[81]
+ wr_data[82] wr_data[83] wr_data[84] wr_data[85] wr_data[86] wr_data[87] wr_data[88]
+ wr_data[89] wr_data[8] wr_data[90] wr_data[91] wr_data[92] wr_data[93] wr_data[94]
+ wr_data[95] wr_data[96] wr_data[97] wr_data[98] wr_data[99] wr_data[9]
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0717__B1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0849__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input127_A wr_data[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input92_A dout0_to_sram[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0613__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0985_ _0638_/X _0984_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1153_/D sky130_fd_sc_hd__mux2_1
Xoutput412 _1082_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[95] sky130_fd_sc_hd__buf_2
Xoutput401 _1072_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[85] sky130_fd_sc_hd__buf_2
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0560__D_N input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0650__A2 _0642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0938__A0 _0938_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0770_ _0777_/A vssd1 vssd1 vccd1 vccd1 _0770_/X sky130_fd_sc_hd__buf_2
XFILLER_5_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1143__GATE_N _0834_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0952__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0968_ _0967_/X _0968_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0968_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _1083_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput264 _1137_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[15] sky130_fd_sc_hd__buf_2
Xoutput253 _0843_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[5] sky130_fd_sc_hd__buf_2
Xoutput275 _1147_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[25] sky130_fd_sc_hd__buf_2
Xoutput286 _1128_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[6] sky130_fd_sc_hd__buf_2
X_0899_ _0898_/X _0899_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0899_/X sky130_fd_sc_hd__mux2_2
Xoutput242 _0851_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[13] sky130_fd_sc_hd__buf_2
Xoutput297 _1093_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[106] sky130_fd_sc_hd__buf_2
XANTENNA__0862__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input194_A wr_data[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A data_to_core_mem[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output309_A _1104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0822_ _1105_/Q _0818_/X input87/X _0819_/X vssd1 vssd1 vccd1 vccd1 _1105_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0753_ _1058_/Q _0749_/X _0801_/B1 _0750_/X vssd1 vssd1 vccd1 vccd1 _1058_/D sky130_fd_sc_hd__a22o_1
X_0684_ _1015_/Q _0679_/X input93/X _0680_/X vssd1 vssd1 vccd1 vccd1 _1015_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_3_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0947__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1098_ _1100_/CLK _1098_/D vssd1 vssd1 vccd1 vccd1 _1098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0857__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input207_A wr_data[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0621__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1021_ _1120_/CLK _1021_/D vssd1 vssd1 vccd1 vccd1 _1021_/Q sky130_fd_sc_hd__dfxtp_1
X_0805_ _0805_/A vssd1 vssd1 vccd1 vccd1 _0805_/X sky130_fd_sc_hd__buf_2
X_0667_ _1002_/Q _0665_/X input79/X _0666_/X vssd1 vssd1 vccd1 vccd1 _1002_/D sky130_fd_sc_hd__a22o_1
X_0736_ _1050_/Q _0707_/A input97/X _0708_/A vssd1 vssd1 vccd1 vccd1 _1050_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0531__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0598_ _0598_/A vssd1 vssd1 vccd1 vccd1 _0598_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input157_A wr_data[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input18_A addr_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0817__A2 _0811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0521_ _0521_/A _0521_/B vssd1 vssd1 vccd1 vccd1 _0522_/C sky130_fd_sc_hd__or2_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0753__B2 _0750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1004_ _1107_/CLK _1004_/D vssd1 vssd1 vccd1 vccd1 _1004_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0960__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0808__A2 _0804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0719_ _1037_/Q _0714_/X input82/X _0715_/X vssd1 vssd1 vccd1 vccd1 _1037_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0744__A1 _1051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0870__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0735__B2 _0708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput120 wr_data[109] vssd1 vssd1 vccd1 vccd1 _0910_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput131 wr_data[119] vssd1 vssd1 vccd1 vccd1 _0950_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput186 wr_data[53] vssd1 vssd1 vccd1 vccd1 _0943_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput197 wr_data[63] vssd1 vssd1 vccd1 vccd1 _0983_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput153 wr_data[23] vssd1 vssd1 vccd1 vccd1 _0952_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput175 wr_data[43] vssd1 vssd1 vccd1 vccd1 _0903_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput142 wr_data[13] vssd1 vssd1 vccd1 vccd1 _0912_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput164 wr_data[33] vssd1 vssd1 vccd1 vccd1 _0863_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__0671__B1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0974__A1 _0974_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0504_ _0507_/A _0507_/C _0501_/A _0503_/A vssd1 vssd1 vccd1 vccd1 _0504_/X sky130_fd_sc_hd__o22a_1
XANTENNA__0726__B2 _0722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0955__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0662__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0717__A1 _1035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0717__B2 _0715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0865__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1138__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0653__B1 _0799_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input85_A dout0_to_sram[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output339_A _1016_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output241_A _0850_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0984_ _0983_/X _0984_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0984_/X sky130_fd_sc_hd__mux2_1
Xoutput402 _1073_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[86] sky130_fd_sc_hd__buf_2
XFILLER_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput413 _1083_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[96] sky130_fd_sc_hd__buf_2
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input237_A wr_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0874__A0 _0874_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0967_ _0966_/X _0967_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0967_/X sky130_fd_sc_hd__mux2_1
Xoutput276 _1148_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[26] sky130_fd_sc_hd__buf_2
Xoutput254 _0844_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[6] sky130_fd_sc_hd__buf_2
Xoutput265 _1138_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[16] sky130_fd_sc_hd__buf_2
X_0898_ _0898_/A0 _0898_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0898_/X sky130_fd_sc_hd__mux2_1
Xoutput287 _1129_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[7] sky130_fd_sc_hd__buf_2
Xoutput243 _0852_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[14] sky130_fd_sc_hd__buf_2
Xoutput298 _1094_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[107] sky130_fd_sc_hd__buf_2
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input187_A wr_data[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input48_A data_to_core_mem[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0619__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0847__A0 _0530_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0821_ _1104_/Q _0818_/X input86/X _0819_/X vssd1 vssd1 vccd1 vccd1 _1104_/D sky130_fd_sc_hd__a22o_1
X_0752_ _1057_/Q _0749_/X _0800_/B1 _0750_/X vssd1 vssd1 vccd1 vccd1 _1057_/D sky130_fd_sc_hd__a22o_1
X_0683_ _1014_/Q _0679_/X input92/X _0680_/X vssd1 vssd1 vccd1 vccd1 _1014_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0963__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1097_ _1114_/CLK _1097_/D vssd1 vssd1 vccd1 vccd1 _1097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0873__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input102_A dout0_to_sram[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0829__B1 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _1116_/CLK sky130_fd_sc_hd__clkbuf_2
X_1020_ _1109_/CLK _1020_/D vssd1 vssd1 vccd1 vccd1 _1020_/Q sky130_fd_sc_hd__dfxtp_1
X_0735_ _1049_/Q _0707_/A input96/X _0708_/A vssd1 vssd1 vccd1 vccd1 _1049_/D sky130_fd_sc_hd__a22o_1
X_0804_ _0804_/A vssd1 vssd1 vccd1 vccd1 _0804_/X sky130_fd_sc_hd__buf_2
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0666_ _0680_/A vssd1 vssd1 vccd1 vccd1 _0666_/X sky130_fd_sc_hd__buf_2
X_0597_ _0857_/S _0597_/B vssd1 vssd1 vccd1 vccd1 _0598_/A sky130_fd_sc_hd__and2_1
XANTENNA__0958__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1149_ _1149_/D _0834_/Y vssd1 vssd1 vccd1 vccd1 _1149_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0868__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0520_ _0521_/A _0517_/A _0521_/B vssd1 vssd1 vccd1 vccd1 _0520_/X sky130_fd_sc_hd__o21a_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0753__A2 _0749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ _1110_/CLK _1003_/D vssd1 vssd1 vccd1 vccd1 _1003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0718_ _1036_/Q _0714_/X input81/X _0715_/X vssd1 vssd1 vccd1 vccd1 _1036_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0649_ _0990_/Q _0642_/X input98/X _0645_/X vssd1 vssd1 vccd1 vccd1 _0990_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1134__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput110 wr_data[0] vssd1 vssd1 vccd1 vccd1 _0860_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0735__A2 _0707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput154 wr_data[24] vssd1 vssd1 vccd1 vccd1 _0956_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput187 wr_data[54] vssd1 vssd1 vccd1 vccd1 _0947_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0627__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput198 wr_data[64] vssd1 vssd1 vccd1 vccd1 _0858_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput176 wr_data[44] vssd1 vssd1 vccd1 vccd1 _0907_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput143 wr_data[14] vssd1 vssd1 vccd1 vccd1 _0916_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input30_A addr_to_core_mem[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput121 wr_data[10] vssd1 vssd1 vccd1 vccd1 _0900_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput132 wr_data[11] vssd1 vssd1 vccd1 vccd1 _0904_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput165 wr_data[34] vssd1 vssd1 vccd1 vccd1 _0867_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0671__B2 _0666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0726__A2 _0721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0503_ _0503_/A vssd1 vssd1 vccd1 vccd1 _0507_/C sky130_fd_sc_hd__inv_2
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0971__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0662__B2 _0659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0717__A2 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0881__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0653__B2 _0652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input78_A dout0_to_sram[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0983_ _0982_/X _0983_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0983_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput414 _1084_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[97] sky130_fd_sc_hd__buf_2
Xoutput403 _1074_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[87] sky130_fd_sc_hd__buf_2
XANTENNA__0883__A1 _0883_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0966__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0876__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input132_A wr_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0562__B1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0966_ _0966_/A0 _0966_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0966_/X sky130_fd_sc_hd__mux2_1
X_0897_ _0594_/X _0896_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1131_/D sky130_fd_sc_hd__mux2_1
Xoutput277 _1149_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[27] sky130_fd_sc_hd__buf_2
Xoutput244 _0853_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[15] sky130_fd_sc_hd__buf_2
Xoutput288 _1130_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[8] sky130_fd_sc_hd__buf_2
Xoutput255 _0845_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[7] sky130_fd_sc_hd__buf_2
Xoutput299 _1095_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[108] sky130_fd_sc_hd__buf_2
Xoutput266 _1139_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[17] sky130_fd_sc_hd__buf_2
XANTENNA__0856__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0792__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0635__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0751_ _1056_/Q _0749_/X _0799_/B1 _0750_/X vssd1 vssd1 vccd1 vccd1 _1056_/D sky130_fd_sc_hd__a22o_1
X_0820_ _1103_/Q _0818_/X input85/X _0819_/X vssd1 vssd1 vccd1 vccd1 _1103_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0783__B1 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0682_ _1013_/Q _0679_/X input91/X _0680_/X vssd1 vssd1 vccd1 vccd1 _1013_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1096_ _1110_/CLK _1096_/D vssd1 vssd1 vccd1 vccd1 _1096_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0838__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0949_ _0620_/X _0948_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1144_/D sky130_fd_sc_hd__mux2_1
XANTENNA__0774__B1 input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0829__B2 _0826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0765__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input60_A data_to_core_mem[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1129__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0803_ _1092_/Q _0797_/X _0803_/B1 _0798_/X vssd1 vssd1 vccd1 vccd1 _1092_/D sky130_fd_sc_hd__a22o_1
X_0734_ _1048_/Q _0728_/X input94/X _0729_/X vssd1 vssd1 vccd1 vccd1 _1048_/D sky130_fd_sc_hd__a22o_1
X_0665_ _0679_/A vssd1 vssd1 vccd1 vccd1 _0665_/X sky130_fd_sc_hd__buf_2
X_0596_ _0596_/A vssd1 vssd1 vccd1 vccd1 _0596_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1148_ _1148_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1148_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1079_ _1110_/CLK _1079_/D vssd1 vssd1 vccd1 vccd1 _1079_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0974__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0747__B1 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0884__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1130__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input212_A wr_data[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ _1107_/CLK _1002_/D vssd1 vssd1 vccd1 vccd1 _1002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0969__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0648_ _0989_/Q _0642_/X input95/X _0645_/X vssd1 vssd1 vccd1 vccd1 _0989_/D sky130_fd_sc_hd__a22o_1
X_0717_ _1035_/Q _0714_/X input80/X _0715_/X vssd1 vssd1 vccd1 vccd1 _1035_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0579_ _0857_/S _0579_/B vssd1 vssd1 vccd1 vccd1 _0580_/A sky130_fd_sc_hd__and2_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0879__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _1120_/CLK sky130_fd_sc_hd__clkbuf_2
Xinput133 wr_data[120] vssd1 vssd1 vccd1 vccd1 _0954_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput122 wr_data[110] vssd1 vssd1 vccd1 vccd1 _0914_/A0 sky130_fd_sc_hd__buf_2
Xinput111 wr_data[100] vssd1 vssd1 vccd1 vccd1 _0874_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput144 wr_data[15] vssd1 vssd1 vccd1 vccd1 _0920_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput100 dout0_to_sram[5] vssd1 vssd1 vccd1 vccd1 _0799_/B1 sky130_fd_sc_hd__buf_4
XANTENNA_input162_A wr_data[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput177 wr_data[45] vssd1 vssd1 vccd1 vccd1 _0911_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput155 wr_data[25] vssd1 vssd1 vccd1 vccd1 _0960_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input23_A addr_to_core_mem[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput188 wr_data[55] vssd1 vssd1 vccd1 vccd1 _0951_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput166 wr_data[35] vssd1 vssd1 vccd1 vccd1 _0871_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput199 wr_data[65] vssd1 vssd1 vccd1 vccd1 _0862_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0671__A2 _0665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0502_ _1119_/Q input12/X _0497_/Y _0499_/X vssd1 vssd1 vccd1 vccd1 _0503_/A sky130_fd_sc_hd__a22o_1
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0662__A2 _0658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0653__A2 _0651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0982_ _0982_/A0 _0982_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0982_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput404 _1075_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[88] sky130_fd_sc_hd__buf_2
Xoutput415 _1085_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[98] sky130_fd_sc_hd__buf_2
XANTENNA__0982__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input125_A wr_data[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0892__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input90_A dout0_to_sram[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0562__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output344_A _1020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0965_ _0628_/X _0964_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1148_/D sky130_fd_sc_hd__mux2_1
X_0896_ _0895_/X _0896_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0896_/X sky130_fd_sc_hd__mux2_1
Xoutput289 _1131_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[9] sky130_fd_sc_hd__buf_2
Xoutput245 _0854_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[16] sky130_fd_sc_hd__buf_2
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0977__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput256 _0846_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[8] sky130_fd_sc_hd__buf_2
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput267 _1140_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[18] sky130_fd_sc_hd__buf_2
Xoutput278 _1150_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[28] sky130_fd_sc_hd__buf_2
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0887__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0792__A1 _1083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0792__B2 _0791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1125__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0750_ _0757_/A vssd1 vssd1 vccd1 vccd1 _0750_/X sky130_fd_sc_hd__clkbuf_4
X_0681_ _1012_/Q _0679_/X input90/X _0680_/X vssd1 vssd1 vccd1 vccd1 _1012_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1095_ _1112_/CLK _1095_/D vssd1 vssd1 vccd1 vccd1 _1095_/Q sky130_fd_sc_hd__dfxtp_1
X_0948_ _0947_/X _0948_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0948_/X sky130_fd_sc_hd__mux2_1
X_0879_ _0878_/X _0879_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0879_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0774__B2 _0771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0829__A2 _0825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input192_A wr_data[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input53_A data_to_core_mem[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0802_ _1091_/Q _0797_/X _0802_/B1 _0798_/X vssd1 vssd1 vccd1 vccd1 _1091_/D sky130_fd_sc_hd__a22o_1
X_0733_ _1047_/Q _0728_/X input93/X _0729_/X vssd1 vssd1 vccd1 vccd1 _1047_/D sky130_fd_sc_hd__a22o_1
X_0664_ _1001_/Q _0658_/X input78/X _0659_/X vssd1 vssd1 vccd1 vccd1 _1001_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0595_ _0857_/S _0595_/B vssd1 vssd1 vccd1 vccd1 _0596_/A sky130_fd_sc_hd__and2_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1147_ _1147_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1147_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_1_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1078_ _1112_/CLK _1078_/D vssd1 vssd1 vccd1 vccd1 _1078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input205_A wr_data[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0683__B1 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0674__B1 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1001_ _1110_/CLK _1001_/D vssd1 vssd1 vccd1 vccd1 _1001_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0977__A1 _0976_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0716_ _1034_/Q _0714_/X input79/X _0715_/X vssd1 vssd1 vccd1 vccd1 _1034_/D sky130_fd_sc_hd__a22o_1
X_0647_ _0988_/Q _0642_/X input84/X _0645_/X vssd1 vssd1 vccd1 vccd1 _0988_/D sky130_fd_sc_hd__a22o_1
X_0578_ _0578_/A vssd1 vssd1 vccd1 vccd1 _0578_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0901__A1 _0900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0985__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0968__A1 _0968_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput167 wr_data[36] vssd1 vssd1 vccd1 vccd1 _0875_/A1 sky130_fd_sc_hd__buf_2
Xinput178 wr_data[46] vssd1 vssd1 vccd1 vccd1 _0915_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput123 wr_data[111] vssd1 vssd1 vccd1 vccd1 _0918_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput156 wr_data[26] vssd1 vssd1 vccd1 vccd1 _0964_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput112 wr_data[101] vssd1 vssd1 vccd1 vccd1 _0878_/A0 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input155_A wr_data[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0895__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput101 dout0_to_sram[6] vssd1 vssd1 vccd1 vccd1 _0800_/B1 sky130_fd_sc_hd__clkbuf_4
Xinput145 wr_data[16] vssd1 vssd1 vccd1 vccd1 _0924_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput134 wr_data[121] vssd1 vssd1 vccd1 vccd1 _0958_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput189 wr_data[56] vssd1 vssd1 vccd1 vccd1 _0955_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0656__B1 _0802_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_A addr_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output374_A _1047_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0501_ _0501_/A vssd1 vssd1 vccd1 vccd1 _0507_/A sky130_fd_sc_hd__inv_2
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0647__B1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_A addr_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0810__B1 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0981_ _0636_/X _0980_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1152_/D sky130_fd_sc_hd__mux2_1
XANTENNA__0801__B1 _0801_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput405 _1076_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[89] sky130_fd_sc_hd__buf_2
Xoutput416 _1086_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[99] sky130_fd_sc_hd__buf_2
XFILLER_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input118_A wr_data[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input83_A dout0_to_sram[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0562__A2 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1121__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0964_ _0963_/X _0964_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0964_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput246 _0855_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[17] sky130_fd_sc_hd__buf_2
Xoutput268 _1141_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[19] sky130_fd_sc_hd__buf_2
X_0895_ _0894_/X _0895_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0895_/X sky130_fd_sc_hd__mux2_1
Xoutput257 _0847_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[9] sky130_fd_sc_hd__buf_2
Xoutput279 _1151_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[29] sky130_fd_sc_hd__buf_2
XFILLER_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0792__A2 _0788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input235_A wr_data[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0680_ _0680_/A vssd1 vssd1 vccd1 vccd1 _0680_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1094_ _1094_/CLK _1094_/D vssd1 vssd1 vccd1 vccd1 _1094_/Q sky130_fd_sc_hd__dfxtp_1
X_0947_ _0946_/X _0947_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0947_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0878_ _0878_/A0 _0878_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0878_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0774__A2 _0770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0898__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input185_A wr_data[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input46_A data_to_core_mem[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0801_ _1090_/Q _0797_/X _0801_/B1 _0798_/X vssd1 vssd1 vccd1 vccd1 _1090_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0663_ _1000_/Q _0658_/X input77/X _0659_/X vssd1 vssd1 vccd1 vccd1 _1000_/D sky130_fd_sc_hd__a22o_1
X_0732_ _1046_/Q _0728_/X input92/X _0729_/X vssd1 vssd1 vccd1 vccd1 _1046_/D sky130_fd_sc_hd__a22o_1
X_0594_ _0594_/A vssd1 vssd1 vccd1 vccd1 _0594_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1146_ _1146_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1146_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1077_ _1112_/CLK _1077_/D vssd1 vssd1 vccd1 vccd1 _1077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0834__B1_N _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input100_A dout0_to_sram[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1000_ _1114_/CLK _1000_/D vssd1 vssd1 vccd1 vccd1 _1000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0674__B2 _0673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0715_ _0729_/A vssd1 vssd1 vccd1 vccd1 _0715_/X sky130_fd_sc_hd__buf_2
XFILLER_30_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0646_ _0987_/Q _0642_/X input73/X _0645_/X vssd1 vssd1 vccd1 vccd1 _0987_/D sky130_fd_sc_hd__a22o_1
X_0577_ _0857_/S _0577_/B vssd1 vssd1 vccd1 vccd1 _0578_/A sky130_fd_sc_hd__and2_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1129_ _1129_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1129_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput146 wr_data[17] vssd1 vssd1 vccd1 vccd1 _0928_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput102 dout0_to_sram[7] vssd1 vssd1 vccd1 vccd1 _0801_/B1 sky130_fd_sc_hd__buf_4
Xinput113 wr_data[102] vssd1 vssd1 vccd1 vccd1 _0882_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput135 wr_data[122] vssd1 vssd1 vccd1 vccd1 _0962_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput168 wr_data[37] vssd1 vssd1 vccd1 vccd1 _0879_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput124 wr_data[112] vssd1 vssd1 vccd1 vccd1 _0922_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput179 wr_data[47] vssd1 vssd1 vccd1 vccd1 _0919_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput157 wr_data[27] vssd1 vssd1 vccd1 vccd1 _0968_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input148_A wr_data[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0656__B2 _0652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0500_ _0497_/Y _0499_/X _0497_/Y _0499_/X vssd1 vssd1 vccd1 vccd1 _0500_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__0647__B2 _0645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0895__A1 _0895_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0886__A1 _0886_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0629_ _0857_/S _0629_/B vssd1 vssd1 vccd1 vccd1 _0630_/A sky130_fd_sc_hd__and2_1
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0810__B2 _0805_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0980_ _0979_/X _0980_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0980_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput406 _0995_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[8] sky130_fd_sc_hd__buf_2
Xoutput417 _0996_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0556__B1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0859__A1 _0859_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0795__B1 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input76_A dout0_to_sram[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0963_ _0962_/X _0963_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0963_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0894_ _0894_/A0 _0894_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0894_/X sky130_fd_sc_hd__mux2_1
Xoutput258 _1122_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[0] sky130_fd_sc_hd__buf_2
Xoutput269 _1123_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[1] sky130_fd_sc_hd__buf_2
Xoutput247 _0856_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[18] sky130_fd_sc_hd__buf_2
XANTENNA__0710__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input130_A wr_data[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input228_A wr_data[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0768__B1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1093_ _1094_/CLK _1093_/D vssd1 vssd1 vccd1 vccd1 _1093_/Q sky130_fd_sc_hd__dfxtp_1
X_0946_ _0946_/A0 _0946_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0946_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0759__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0877_ _0584_/X _0876_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1126_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input178_A wr_data[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0922__A0 _0922_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A addr_to_core_mem[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0800_ _1089_/Q _0797_/X _0800_/B1 _0798_/X vssd1 vssd1 vccd1 vccd1 _1089_/D sky130_fd_sc_hd__a22o_1
X_0731_ _1045_/Q _0728_/X input91/X _0729_/X vssd1 vssd1 vccd1 vccd1 _1045_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0662_ _0999_/Q _0658_/X input76/X _0659_/X vssd1 vssd1 vccd1 vccd1 _0999_/D sky130_fd_sc_hd__a22o_1
X_0593_ _0857_/S _0593_/B vssd1 vssd1 vccd1 vccd1 _0594_/A sky130_fd_sc_hd__and2_1
X_1145_ _1145_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1145_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1076_ _1094_/CLK _1076_/D vssd1 vssd1 vccd1 vccd1 _1076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0929_ _0610_/X _0928_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1139_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output312_A _0998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0674__A2 _0672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0645_ _0659_/A vssd1 vssd1 vccd1 vccd1 _0645_/X sky130_fd_sc_hd__buf_2
X_0714_ _0728_/A vssd1 vssd1 vccd1 vccd1 _0714_/X sky130_fd_sc_hd__buf_2
X_0576_ _0576_/A vssd1 vssd1 vccd1 vccd1 _0982_/S sky130_fd_sc_hd__buf_12
XFILLER_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1128_ _1128_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1128_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0583__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1059_ _1112_/CLK _1059_/D vssd1 vssd1 vccd1 vccd1 _1059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput103 dout0_to_sram[8] vssd1 vssd1 vccd1 vccd1 _0802_/B1 sky130_fd_sc_hd__buf_6
Xinput169 wr_data[38] vssd1 vssd1 vccd1 vccd1 _0883_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput158 wr_data[28] vssd1 vssd1 vccd1 vccd1 _0972_/A1 sky130_fd_sc_hd__buf_2
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput136 wr_data[123] vssd1 vssd1 vccd1 vccd1 _0966_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput114 wr_data[103] vssd1 vssd1 vccd1 vccd1 _0886_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput147 wr_data[18] vssd1 vssd1 vccd1 vccd1 _0932_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput125 wr_data[113] vssd1 vssd1 vccd1 vccd1 _0926_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input210_A wr_data[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0656__A2 _0651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0647__A2 _0642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0628_ _0628_/A vssd1 vssd1 vccd1 vccd1 _0628_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0559_ input8/X input9/X _0554_/A _0558_/X vssd1 vssd1 vccd1 vccd1 _0559_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0810__A2 _0804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input160_A wr_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A addr_to_core_mem[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0568__A_N _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput418 _0986_/S vssd1 vssd1 vccd1 vccd1 ready sky130_fd_sc_hd__buf_2
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput407 _1077_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[90] sky130_fd_sc_hd__buf_2
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0795__A1 _1086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0795__B2 _0791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input69_A data_to_core_mem[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0962_ _0962_/A0 _0962_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0962_/X sky130_fd_sc_hd__mux2_1
X_0893_ _0592_/X _0892_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1130_/D sky130_fd_sc_hd__mux2_2
Xoutput259 _1132_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[10] sky130_fd_sc_hd__buf_2
Xoutput248 _0857_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[19] sky130_fd_sc_hd__buf_2
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0710__A1 _1030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0710__B2 _0708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0591__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input123_A wr_data[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1092_ _1107_/CLK _1092_/D vssd1 vssd1 vccd1 vccd1 _1092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0945_ _0618_/X _0944_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1143_/D sky130_fd_sc_hd__mux2_1
X_0876_ _0875_/X _0876_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0876_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0695__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0922__A1 _0922_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0686__B1 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0730_ _1044_/Q _0728_/X input90/X _0729_/X vssd1 vssd1 vccd1 vccd1 _1044_/D sky130_fd_sc_hd__a22o_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0661_ _0998_/Q _0658_/X input75/X _0659_/X vssd1 vssd1 vccd1 vccd1 _0998_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0592_ _0592_/A vssd1 vssd1 vccd1 vccd1 _0592_/X sky130_fd_sc_hd__clkbuf_1
X_1075_ _1075_/CLK _1075_/D vssd1 vssd1 vccd1 vccd1 _1075_/Q sky130_fd_sc_hd__dfxtp_1
X_1144_ _1144_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1144_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0677__B1 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0859_ _0858_/X _0859_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0859_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0928_ _0927_/X _0928_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0928_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0668__B1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input190_A wr_data[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input51_A data_to_core_mem[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0831__B1 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0644_ _0680_/A vssd1 vssd1 vccd1 vccd1 _0659_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0713_ _1033_/Q _0707_/X input78/X _0708_/X vssd1 vssd1 vccd1 vccd1 _1033_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0575_ _0575_/A _0575_/B _1119_/Q _0575_/D vssd1 vssd1 vccd1 vccd1 _0576_/A sky130_fd_sc_hd__and4_1
X_1127_ _1127_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1127_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1058_ _1114_/CLK _1058_/D vssd1 vssd1 vccd1 vccd1 _1058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0822__B1 input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput126 wr_data[114] vssd1 vssd1 vccd1 vccd1 _0930_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput115 wr_data[104] vssd1 vssd1 vccd1 vccd1 _0890_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput104 dout0_to_sram[9] vssd1 vssd1 vccd1 vccd1 _0803_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput137 wr_data[124] vssd1 vssd1 vccd1 vccd1 _0970_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput148 wr_data[19] vssd1 vssd1 vccd1 vccd1 _0936_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput159 wr_data[29] vssd1 vssd1 vccd1 vccd1 _0976_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0813__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input203_A wr_data[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input99_A dout0_to_sram[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output255_A _0845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0627_ _0857_/S _0627_/B vssd1 vssd1 vccd1 vccd1 _0628_/A sky130_fd_sc_hd__and2_1
X_0558_ _0560_/A _0560_/C _0560_/B vssd1 vssd1 vccd1 vccd1 _0558_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0489_ _0488_/Y _0986_/S _0487_/A _0487_/B vssd1 vssd1 vccd1 vccd1 _0492_/A sky130_fd_sc_hd__a211o_1
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input153_A wr_data[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A addr_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput408 _1078_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[91] sky130_fd_sc_hd__buf_2
Xoutput419 _1121_/Q vssd1 vssd1 vccd1 vccd1 we_to_sram sky130_fd_sc_hd__buf_2
XFILLER_35_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0589__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_A addr_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0795__A2 _0788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0961_ _0626_/X _0960_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1147_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0901__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0892_ _0891_/X _0892_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0892_/X sky130_fd_sc_hd__mux2_1
Xoutput249 _0839_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[1] sky130_fd_sc_hd__buf_2
Xoutput238 _0838_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[0] sky130_fd_sc_hd__buf_2
XANTENNA__0710__A2 _0707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A wr_data[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input81_A dout0_to_sram[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1091_ _1091_/CLK _1091_/D vssd1 vssd1 vccd1 vccd1 _1091_/Q sky130_fd_sc_hd__dfxtp_1
X_0944_ _0943_/X _0944_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0944_/X sky130_fd_sc_hd__mux2_1
X_0875_ _0874_/X _0875_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0875_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0695__A1 _1019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input233_A wr_data[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0686__A1 _1017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0591_ _0857_/S _0591_/B vssd1 vssd1 vccd1 vccd1 _0592_/A sky130_fd_sc_hd__and2_1
X_0660_ _0997_/Q _0658_/X input74/X _0659_/X vssd1 vssd1 vccd1 vccd1 _0997_/D sky130_fd_sc_hd__a22o_1
X_1143_ _1143_/D _0834_/Y vssd1 vssd1 vccd1 vccd1 _1143_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1074_ _1075_/CLK _1074_/D vssd1 vssd1 vccd1 vccd1 _1074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0677__B2 _0673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0677__A1 _1010_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0927_ _0926_/X _0927_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0927_/X sky130_fd_sc_hd__mux2_1
X_0858_ _0858_/A0 _0858_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0858_/X sky130_fd_sc_hd__mux2_1
X_0789_ _0825_/A vssd1 vssd1 vccd1 vccd1 _0826_/A sky130_fd_sc_hd__inv_2
XANTENNA__0597__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0668__B2 _0666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input183_A wr_data[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input44_A data_to_core_mem[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0831__B2 _0826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0643_ _0679_/A vssd1 vssd1 vccd1 vccd1 _0680_/A sky130_fd_sc_hd__inv_2
X_0712_ _1032_/Q _0707_/X input77/X _0708_/X vssd1 vssd1 vccd1 vccd1 _1032_/D sky130_fd_sc_hd__a22o_1
X_0574_ _0574_/A vssd1 vssd1 vccd1 vccd1 _0983_/S sky130_fd_sc_hd__buf_12
XFILLER_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1126_ _1126_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1126_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0822__B2 _0819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1057_ _1111_/CLK _1057_/D vssd1 vssd1 vccd1 vccd1 _1057_/Q sky130_fd_sc_hd__dfxtp_1
Xinput116 wr_data[105] vssd1 vssd1 vccd1 vccd1 _0894_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput105 is_loading_memory_into_core vssd1 vssd1 vccd1 vccd1 _0857_/S sky130_fd_sc_hd__buf_12
Xinput127 wr_data[115] vssd1 vssd1 vccd1 vccd1 _0934_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput149 wr_data[1] vssd1 vssd1 vccd1 vccd1 _0864_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput138 wr_data[125] vssd1 vssd1 vccd1 vccd1 _0974_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0813__B2 _0812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1151__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output248_A _0857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0904__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0557_ input9/X vssd1 vssd1 vccd1 vccd1 _0560_/B sky130_fd_sc_hd__inv_2
X_0626_ _0626_/A vssd1 vssd1 vccd1 vccd1 _0626_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1109_ _1109_/CLK _1109_/D vssd1 vssd1 vccd1 vccd1 _1109_/Q sky130_fd_sc_hd__dfxtp_1
X_0488_ _0568_/C vssd1 vssd1 vccd1 vccd1 _0488_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input146_A wr_data[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0731__B1 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput409 _1079_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[92] sky130_fd_sc_hd__buf_2
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0713__B1 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0609_ _0857_/S _0609_/B vssd1 vssd1 vccd1 vccd1 _0610_/A sky130_fd_sc_hd__and2_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0704__B1 _0801_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0960_ _0959_/X _0960_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0960_/X sky130_fd_sc_hd__mux2_1
Xoutput239 _0848_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[10] sky130_fd_sc_hd__buf_2
X_0891_ _0890_/X _0891_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0891_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input74_A dout0_to_sram[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1090_ _1091_/CLK _1090_/D vssd1 vssd1 vccd1 vccd1 _1090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0943_ _0942_/X _0943_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0943_/X sky130_fd_sc_hd__mux2_1
X_0874_ _0874_/A0 _0874_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0874_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0912__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0907__A0 _0906_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input226_A wr_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0590_ _0590_/A vssd1 vssd1 vccd1 vccd1 _0590_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1142_ _1142_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1142_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_1_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0677__A2 _0672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1073_ _1091_/CLK _1073_/D vssd1 vssd1 vccd1 vccd1 _1073_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0907__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0857_ _0565_/X input31/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0857_/X sky130_fd_sc_hd__mux2_2
X_0926_ _0926_/A0 _0926_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0926_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1146__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0788_ _0804_/A vssd1 vssd1 vccd1 vccd1 _0788_/X sky130_fd_sc_hd__buf_2
XFILLER_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0597__B _0597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0668__A2 _0665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input176_A wr_data[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input37_A addr_to_core_mem[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0711_ _1031_/Q _0707_/X input76/X _0708_/X vssd1 vssd1 vccd1 vccd1 _1031_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0831__A2 _0825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0642_ _0658_/A vssd1 vssd1 vccd1 vccd1 _0642_/X sky130_fd_sc_hd__buf_2
X_0573_ _0575_/A _0575_/B _1119_/Q _1117_/Q vssd1 vssd1 vccd1 vccd1 _0574_/A sky130_fd_sc_hd__and4_1
X_1125_ _1125_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1125_/Q sky130_fd_sc_hd__dlxtn_1
X_1056_ _1109_/CLK _1056_/D vssd1 vssd1 vccd1 vccd1 _1056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0909_ _0600_/X _0908_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1134_/D sky130_fd_sc_hd__mux2_1
Xinput128 wr_data[116] vssd1 vssd1 vccd1 vccd1 _0938_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput106 requested vssd1 vssd1 vccd1 vccd1 _0568_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput139 wr_data[126] vssd1 vssd1 vccd1 vccd1 _0978_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput117 wr_data[106] vssd1 vssd1 vccd1 vccd1 _0898_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0813__A2 _0811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0920__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0625_ _0857_/S _0625_/B vssd1 vssd1 vccd1 vccd1 _0626_/A sky130_fd_sc_hd__and2_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0556_ _0560_/A _0560_/C input8/X _0554_/A vssd1 vssd1 vccd1 vccd1 _0556_/X sky130_fd_sc_hd__o22a_1
X_0487_ _0487_/A _0487_/B _0487_/C vssd1 vssd1 vccd1 vccd1 _1119_/D sky130_fd_sc_hd__nor3_1
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1039_ _1100_/CLK _1039_/D vssd1 vssd1 vccd1 vccd1 _1039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1108_ _1111_/CLK _1108_/D vssd1 vssd1 vccd1 vccd1 _1108_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0559__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input139_A wr_data[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0970__A1 _0970_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0915__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0608_ _0608_/A vssd1 vssd1 vccd1 vccd1 _0608_/X sky130_fd_sc_hd__clkbuf_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0539_ _0539_/A vssd1 vssd1 vccd1 vccd1 _0539_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0713__B2 _0708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0952__A1 _0952_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0890_ _0890_/A0 _0890_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0890_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0698__B1 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input67_A data_to_core_mem[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0861__A0 _0567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0942_ _0942_/A0 _0942_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0942_/X sky130_fd_sc_hd__mux2_1
X_0873_ _0582_/X _0872_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1125_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1142__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0852__A0 _0548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input219_A wr_data[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input121_A wr_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1141_ _1141_/D _0834_/Y vssd1 vssd1 vccd1 vccd1 _1141_/Q sky130_fd_sc_hd__dlxtn_1
X_1072_ _1075_/CLK _1072_/D vssd1 vssd1 vccd1 vccd1 _1072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0923__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0856_ _0563_/Y input30/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0856_/X sky130_fd_sc_hd__mux2_2
X_0787_ _0825_/A vssd1 vssd1 vccd1 vccd1 _0804_/A sky130_fd_sc_hd__clkbuf_2
X_0925_ _0608_/X _0924_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1138_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input169_A wr_data[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput390 _1062_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[75] sky130_fd_sc_hd__buf_2
XFILLER_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0816__B1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0641_ _0679_/A vssd1 vssd1 vccd1 vccd1 _0658_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0710_ _1030_/Q _0707_/X input75/X _0708_/X vssd1 vssd1 vccd1 vccd1 _1030_/D sky130_fd_sc_hd__a22o_1
X_0572_ _0572_/A vssd1 vssd1 vccd1 vccd1 _0984_/S sky130_fd_sc_hd__buf_12
XANTENNA__0918__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1055_ _1083_/CLK _1055_/D vssd1 vssd1 vccd1 vccd1 _1055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1124_ _1124_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1124_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0807__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0908_ _0907_/X _0908_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0908_/X sky130_fd_sc_hd__mux2_1
X_0839_ _0500_/X input32/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0839_/X sky130_fd_sc_hd__mux2_4
Xinput118 wr_data[107] vssd1 vssd1 vccd1 vccd1 _0902_/A0 sky130_fd_sc_hd__buf_2
XFILLER_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput107 reset vssd1 vssd1 vccd1 vccd1 _0487_/B sky130_fd_sc_hd__clkbuf_2
Xinput129 wr_data[117] vssd1 vssd1 vccd1 vccd1 _0942_/A0 sky130_fd_sc_hd__clkbuf_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0624_ _0624_/A vssd1 vssd1 vccd1 vccd1 _0624_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0555_ input8/X vssd1 vssd1 vccd1 vccd1 _0560_/A sky130_fd_sc_hd__inv_2
X_0486_ _1119_/Q _1117_/Q _0571_/C _0484_/B vssd1 vssd1 vccd1 vccd1 _0487_/C sky130_fd_sc_hd__a22oi_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1107_ _1107_/CLK _1107_/D vssd1 vssd1 vccd1 vccd1 _1107_/Q sky130_fd_sc_hd__dfxtp_1
X_1038_ _1083_/CLK _1038_/D vssd1 vssd1 vccd1 vccd1 _1038_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0559__A2 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input97_A dout0_to_sram[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input201_A wr_data[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0931__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0538_ _0535_/X _0551_/D vssd1 vssd1 vccd1 vccd1 _0539_/A sky130_fd_sc_hd__and2b_1
X_0607_ _0857_/S _0607_/B vssd1 vssd1 vccd1 vccd1 _0608_/A sky130_fd_sc_hd__and2_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0713__A2 _0707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0841__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1137__GATE_N _0834_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input151_A wr_data[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1123__D _1123_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A addr_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0926__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_A addr_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0870__A1 _0870_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input199_A wr_data[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0941_ _0616_/X _0940_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1142_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0872_ _0871_/X _0872_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0872_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0510__A _0510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input114_A wr_data[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output333_A _1010_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1071_ _1091_/CLK _1071_/D vssd1 vssd1 vccd1 vccd1 _1071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1140_ _1140_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1140_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_1_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0924_ _0923_/X _0924_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0924_/X sky130_fd_sc_hd__mux2_1
X_0855_ _0559_/Y input29/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0855_/X sky130_fd_sc_hd__mux2_1
X_0786_ _0786_/A _0786_/B vssd1 vssd1 vccd1 vccd1 _0825_/A sky130_fd_sc_hd__or2_2
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput391 _1063_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[76] sky130_fd_sc_hd__buf_2
Xoutput380 _1053_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[66] sky130_fd_sc_hd__buf_2
XANTENNA__0761__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input231_A wr_data[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0816__B2 _0812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1131__D _1131_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0640_ _1115_/Q _1116_/Q vssd1 vssd1 vccd1 vccd1 _0679_/A sky130_fd_sc_hd__or2_1
X_0571_ _0575_/A _1118_/Q _0571_/C vssd1 vssd1 vccd1 vccd1 _0572_/A sky130_fd_sc_hd__and3_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0752__B1 _0800_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0934__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1123_ _1123_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1123_/Q sky130_fd_sc_hd__dlxtn_1
X_1054_ _1116_/CLK _1054_/D vssd1 vssd1 vccd1 vccd1 _1054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0807__B2 _0805_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0807__A1 _1094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0907_ _0906_/X _0907_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0907_/X sky130_fd_sc_hd__mux2_1
Xinput108 reset_mem_req vssd1 vssd1 vccd1 vccd1 _0487_/A sky130_fd_sc_hd__clkbuf_4
X_0769_ _1070_/Q _0763_/X input83/X _0764_/X vssd1 vssd1 vccd1 vccd1 _1070_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0838_ _0498_/Y input21/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0838_/X sky130_fd_sc_hd__mux2_2
XFILLER_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput119 wr_data[108] vssd1 vssd1 vccd1 vccd1 _0906_/A0 sky130_fd_sc_hd__clkbuf_1
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0844__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0982__A0 _0982_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input181_A wr_data[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input42_A data_to_core_mem[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0734__B1 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0623_ _0857_/S _0623_/B vssd1 vssd1 vccd1 vccd1 _0624_/A sky130_fd_sc_hd__and2_1
X_0554_ _0554_/A _0554_/B vssd1 vssd1 vccd1 vccd1 _0554_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__0725__B1 input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0485_ _0485_/A vssd1 vssd1 vccd1 vccd1 _0571_/C sky130_fd_sc_hd__inv_2
XANTENNA__0929__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0489__C1 _0487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1106_ _1106_/CLK _1106_/D vssd1 vssd1 vccd1 vccd1 _1106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1037_ _1107_/CLK _1037_/D vssd1 vssd1 vccd1 vccd1 _1037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 dout0_to_sram[25] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0716__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0839__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1133__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0603__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output413_A _1083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0513__A _0513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0606_ _0606_/A vssd1 vssd1 vccd1 vccd1 _0606_/X sky130_fd_sc_hd__clkbuf_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0537_ _0537_/A _0537_/B _0537_/C _0537_/D vssd1 vssd1 vccd1 vccd1 _0551_/D sky130_fd_sc_hd__or4_2
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input144_A wr_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0942__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0852__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0940_ _0939_/X _0940_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0940_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0871_ _0870_/X _0871_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0871_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0937__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0701__A _0708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0847__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input107_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1129__D _1129_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0611__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input72_A data_to_core_mem[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1070_ _1106_/CLK _1070_/D vssd1 vssd1 vccd1 vccd1 _1070_/Q sky130_fd_sc_hd__dfxtp_1
X_0854_ _0556_/X input28/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0854_/X sky130_fd_sc_hd__mux2_1
X_0923_ _0922_/X _0923_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0923_/X sky130_fd_sc_hd__mux2_2
X_0785_ _1082_/Q _0756_/A input97/X _0757_/A vssd1 vssd1 vccd1 vccd1 _1082_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput392 _1064_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[77] sky130_fd_sc_hd__buf_2
Xoutput370 _1044_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[57] sky130_fd_sc_hd__buf_2
Xoutput381 _1054_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[67] sky130_fd_sc_hd__buf_2
XFILLER_10_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0816__A2 _0811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input224_A wr_data[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1128__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0570_ _1120_/Q vssd1 vssd1 vccd1 vccd1 _0575_/A sky130_fd_sc_hd__inv_2
X_1122_ _1122_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1122_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0752__B2 _0750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1053_ _1075_/CLK _1053_/D vssd1 vssd1 vccd1 vccd1 _1053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0807__A2 _0804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0950__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0906_ _0906_/A0 _0906_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0906_/X sky130_fd_sc_hd__mux2_1
X_0837_ vssd1 vssd1 vccd1 vccd1 _0837_/HI spare_wen0_to_sram sky130_fd_sc_hd__conb_1
Xinput109 we vssd1 vssd1 vccd1 vccd1 _0568_/B sky130_fd_sc_hd__clkbuf_2
X_0768_ _1069_/Q _0763_/X input82/X _0764_/X vssd1 vssd1 vccd1 vccd1 _1069_/D sky130_fd_sc_hd__a22o_1
X_0699_ _1023_/Q _0691_/X input99/X _0694_/X vssd1 vssd1 vccd1 vccd1 _1023_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0860__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input174_A wr_data[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input35_A addr_to_core_mem[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0670__B1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0622_ _0622_/A vssd1 vssd1 vccd1 vccd1 _0622_/X sky130_fd_sc_hd__clkbuf_1
X_0553_ _0550_/A _0547_/A _0550_/B vssd1 vssd1 vccd1 vccd1 _0554_/B sky130_fd_sc_hd__o21a_1
XANTENNA__0725__B2 _0722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0484_ _0485_/A _0484_/B vssd1 vssd1 vccd1 vccd1 _0986_/S sky130_fd_sc_hd__nor2_4
XANTENNA__0945__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1105_ _1113_/CLK _1105_/D vssd1 vssd1 vccd1 vccd1 _1105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0489__B1 _0487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1036_ _1106_/CLK _1036_/D vssd1 vssd1 vccd1 vccd1 _1036_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0661__B1 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput91 dout0_to_sram[26] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__buf_4
Xinput80 dout0_to_sram[16] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__buf_2
XANTENNA__0716__B2 _0715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0855__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output239_A _0848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0946__A1 _0946_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0605_ _0857_/S _0605_/B vssd1 vssd1 vccd1 vccd1 _0606_/A sky130_fd_sc_hd__and2_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0536_ _0536_/A _0536_/B vssd1 vssd1 vccd1 vccd1 _0537_/C sky130_fd_sc_hd__or2_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1019_ _1111_/CLK _1019_/D vssd1 vssd1 vccd1 vccd1 _1019_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input137_A wr_data[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0928__A1 _0928_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0919__A1 _0919_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0519_ _0519_/A vssd1 vssd1 vccd1 vccd1 _0521_/B sky130_fd_sc_hd__inv_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0846__A0 _0527_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0609__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0870_ _0870_/A0 _0870_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0870_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0953__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0999_ _1114_/CLK _0999_/D vssd1 vssd1 vccd1 vccd1 _0999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0828__B1 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0863__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input65_A data_to_core_mem[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1124__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output319_A _1113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0853_ _0554_/Y input27/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0853_/X sky130_fd_sc_hd__mux2_1
X_0922_ _0922_/A0 _0922_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0922_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0948__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0784_ _1081_/Q _0756_/A input96/X _0757_/A vssd1 vssd1 vccd1 vccd1 _1081_/D sky130_fd_sc_hd__a22o_1
Xinput1 addr_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput393 _1065_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[78] sky130_fd_sc_hd__buf_2
Xoutput382 _1055_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[68] sky130_fd_sc_hd__buf_2
XANTENNA__0858__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput371 _1045_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[58] sky130_fd_sc_hd__buf_2
Xoutput360 _1035_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[48] sky130_fd_sc_hd__buf_2
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input217_A wr_data[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0752__A2 _0749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1052_ _1116_/CLK _1052_/D vssd1 vssd1 vccd1 vccd1 _1052_/Q sky130_fd_sc_hd__dfxtp_1
X_1121_ _1121_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1121_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0836_ vssd1 vssd1 vccd1 vccd1 _0836_/HI csb0_to_sram sky130_fd_sc_hd__conb_1
X_0767_ _1068_/Q _0763_/X input81/X _0764_/X vssd1 vssd1 vccd1 vccd1 _1068_/D sky130_fd_sc_hd__a22o_1
X_0905_ _0598_/X _0904_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1133_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0698_ _1022_/Q _0691_/X input98/X _0694_/X vssd1 vssd1 vccd1 vccd1 _1022_/D sky130_fd_sc_hd__a22o_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0707__A _0707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input167_A wr_data[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input28_A addr_to_core_mem[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0617__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0670__B2 _0666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0621_ _0857_/S _0621_/B vssd1 vssd1 vccd1 vccd1 _0622_/A sky130_fd_sc_hd__and2_1
XFILLER_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0552_ _0560_/C vssd1 vssd1 vccd1 vccd1 _0554_/A sky130_fd_sc_hd__inv_2
XANTENNA__0725__A2 _0721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0483_ _1120_/Q _1118_/Q vssd1 vssd1 vccd1 vccd1 _0484_/B sky130_fd_sc_hd__or2_1
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1104_ _1113_/CLK _1104_/D vssd1 vssd1 vccd1 vccd1 _1104_/Q sky130_fd_sc_hd__dfxtp_1
X_1035_ _1109_/CLK _1035_/D vssd1 vssd1 vccd1 vccd1 _1035_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0961__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0661__B2 _0659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0661__A1 _0998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput81 dout0_to_sram[17] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_2
XANTENNA__0716__A2 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput70 data_to_core_mem[7] vssd1 vssd1 vccd1 vccd1 _0589_/B sky130_fd_sc_hd__clkbuf_1
Xinput92 dout0_to_sram[27] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__buf_2
X_0819_ _0826_/A vssd1 vssd1 vccd1 vccd1 _0819_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0871__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0604_ _0604_/A vssd1 vssd1 vccd1 vccd1 _0604_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0956__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0535_ _0536_/A _0532_/A _0536_/B vssd1 vssd1 vccd1 vccd1 _0535_/X sky130_fd_sc_hd__o21a_1
XANTENNA__0882__A1 _0882_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1018_ _1113_/CLK _1018_/D vssd1 vssd1 vccd1 vccd1 _1018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0866__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input95_A dout0_to_sram[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0518_ _0521_/A _0517_/A _0516_/A _0517_/Y vssd1 vssd1 vccd1 vccd1 _0518_/X sky130_fd_sc_hd__o22a_1
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0855__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input10_A addr_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0625__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0782__B1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0998_ _1106_/CLK _0998_/D vssd1 vssd1 vccd1 vccd1 _0998_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0773__B1 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A addr_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0828__B2 _0826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input197_A wr_data[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input58_A data_to_core_mem[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0921_ _0606_/X _0920_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1137_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0852_ _0548_/X input26/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0852_/X sky130_fd_sc_hd__mux2_1
X_0783_ _1080_/Q _0777_/X input94/X _0778_/X vssd1 vssd1 vccd1 vccd1 _1080_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0755__B1 _0803_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0964__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput2 addr_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0746__B1 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput361 _1036_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[49] sky130_fd_sc_hd__buf_2
Xoutput350 _1026_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[39] sky130_fd_sc_hd__buf_2
Xoutput383 _1056_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[69] sky130_fd_sc_hd__buf_2
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput372 _1046_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[59] sky130_fd_sc_hd__buf_2
Xoutput394 _1066_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[79] sky130_fd_sc_hd__buf_2
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input112_A wr_data[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0874__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1051_ _1083_/CLK _1051_/D vssd1 vssd1 vccd1 vccd1 _1051_/Q sky130_fd_sc_hd__dfxtp_2
X_1120_ _1120_/CLK _1120_/D vssd1 vssd1 vccd1 vccd1 _1120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0904_ _0903_/X _0904_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0904_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0959__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0835_ _0575_/B _0571_/C _0487_/A _0487_/B _0575_/A vssd1 vssd1 vccd1 vccd1 _1120_/D
+ sky130_fd_sc_hd__a2111oi_1
X_0766_ _1067_/Q _0763_/X input80/X _0764_/X vssd1 vssd1 vccd1 vccd1 _1067_/D sky130_fd_sc_hd__a22o_1
X_0697_ _1021_/Q _0691_/X input95/X _0694_/X vssd1 vssd1 vccd1 vccd1 _1021_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0900__A0 _0899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0719__B1 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0869__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0670__A2 _0665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0633__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0620_ _0620_/A vssd1 vssd1 vccd1 vccd1 _0620_/X sky130_fd_sc_hd__clkbuf_1
X_0551_ _0551_/A _0551_/B _0551_/C _0551_/D vssd1 vssd1 vccd1 vccd1 _0560_/C sky130_fd_sc_hd__or4_2
XFILLER_7_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0489__A2 _0986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0482_ _1119_/Q _1117_/Q vssd1 vssd1 vccd1 vccd1 _0485_/A sky130_fd_sc_hd__or2_2
X_1034_ _1100_/CLK _1034_/D vssd1 vssd1 vccd1 vccd1 _1034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1103_ _1106_/CLK _1103_/D vssd1 vssd1 vccd1 vccd1 _1103_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0543__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0661__A2 _0658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput82 dout0_to_sram[18] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__buf_2
Xinput93 dout0_to_sram[28] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__buf_4
X_0749_ _0756_/A vssd1 vssd1 vccd1 vccd1 _0749_/X sky130_fd_sc_hd__clkbuf_4
X_0818_ _0825_/A vssd1 vssd1 vccd1 vccd1 _0818_/X sky130_fd_sc_hd__clkbuf_2
Xinput71 data_to_core_mem[8] vssd1 vssd1 vccd1 vccd1 _0591_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput60 data_to_core_mem[27] vssd1 vssd1 vccd1 vccd1 _0629_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input40_A addr_to_core_mem[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0534_ input3/X vssd1 vssd1 vccd1 vccd1 _0536_/B sky130_fd_sc_hd__inv_2
X_0603_ _0857_/S _0603_/B vssd1 vssd1 vccd1 vccd1 _0604_/A sky130_fd_sc_hd__and2_1
XFILLER_7_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ _1113_/CLK _1017_/D vssd1 vssd1 vccd1 vccd1 _1017_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__0972__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0882__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input88_A dout0_to_sram[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0517_ _0517_/A vssd1 vssd1 vccd1 vccd1 _0517_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0967__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0877__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input142_A wr_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0782__A1 _1079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0773__B2 _0771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0997_ _1110_/CLK _0997_/D vssd1 vssd1 vccd1 vccd1 _0997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0828__A2 _0825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0920_ _0919_/X _0920_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0920_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0851_ _0545_/X input25/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0851_/X sky130_fd_sc_hd__mux2_2
X_0782_ _1079_/Q _0777_/X input93/X _0778_/X vssd1 vssd1 vccd1 vccd1 _1079_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0755__B2 _0750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput3 addr_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0980__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput340 _0989_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[2] sky130_fd_sc_hd__buf_2
Xoutput351 _0990_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[3] sky130_fd_sc_hd__buf_2
Xoutput395 _0994_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[7] sky130_fd_sc_hd__buf_2
Xoutput373 _0992_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[5] sky130_fd_sc_hd__buf_2
Xoutput384 _0993_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_3_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput362 _0991_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input105_A is_loading_memory_into_core vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0890__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0682__B1 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input70_A data_to_core_mem[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1050_ _1100_/CLK _1050_/D vssd1 vssd1 vccd1 vccd1 _1050_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0903_ _0902_/X _0903_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0903_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0976__A1 _0976_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0834_ _0575_/A _0492_/B _0985_/S vssd1 vssd1 vccd1 vccd1 _0834_/Y sky130_fd_sc_hd__a21boi_4
X_0765_ _1066_/Q _0763_/X input79/X _0764_/X vssd1 vssd1 vccd1 vccd1 _1066_/D sky130_fd_sc_hd__a22o_1
X_0696_ _1020_/Q _0691_/X input84/X _0694_/X vssd1 vssd1 vccd1 vccd1 _1020_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0975__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0664__B1 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0719__B2 _0715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0655__B1 _0801_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0885__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input222_A wr_data[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0958__A1 _0958_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0550_ _0550_/A _0550_/B vssd1 vssd1 vccd1 vccd1 _0551_/C sky130_fd_sc_hd__or2_1
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1102_ _1109_/CLK _1102_/D vssd1 vssd1 vccd1 vccd1 _1102_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0894__A0 _0894_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0646__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1033_ _1109_/CLK _1033_/D vssd1 vssd1 vccd1 vccd1 _1033_/Q sky130_fd_sc_hd__dfxtp_1
Xinput61 data_to_core_mem[28] vssd1 vssd1 vccd1 vccd1 _0631_/B sky130_fd_sc_hd__clkbuf_1
X_0817_ _1102_/Q _0811_/X input83/X _0812_/X vssd1 vssd1 vccd1 vccd1 _1102_/D sky130_fd_sc_hd__a22o_1
Xinput50 data_to_core_mem[18] vssd1 vssd1 vccd1 vccd1 _0611_/B sky130_fd_sc_hd__clkbuf_1
Xinput72 data_to_core_mem[9] vssd1 vssd1 vccd1 vccd1 _0593_/B sky130_fd_sc_hd__clkbuf_1
Xinput83 dout0_to_sram[19] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__buf_2
X_0748_ _1055_/Q _0740_/X input99/X _0743_/X vssd1 vssd1 vccd1 vccd1 _1055_/D sky130_fd_sc_hd__a22o_1
Xinput94 dout0_to_sram[29] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__buf_2
X_0679_ _0679_/A vssd1 vssd1 vccd1 vccd1 _0679_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0885__A0 _0588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input172_A wr_data[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A addr_to_core_mem[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0800__B1 _0800_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0533_ _0536_/A _0532_/A input2/X _0532_/Y vssd1 vssd1 vccd1 vccd1 _0533_/X sky130_fd_sc_hd__o22a_1
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0602_ _0602_/A vssd1 vssd1 vccd1 vccd1 _0602_/X sky130_fd_sc_hd__clkbuf_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0867__A0 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ _1094_/CLK _1016_/D vssd1 vssd1 vccd1 vccd1 _1016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_1_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0516_ _0516_/A vssd1 vssd1 vccd1 vccd1 _0521_/A sky130_fd_sc_hd__inv_2
XANTENNA__0549__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0983__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input135_A wr_data[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0893__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0996_ _1094_/CLK _0996_/D vssd1 vssd1 vccd1 vccd1 _0996_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0773__A2 _0770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0978__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0888__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0850_ _0542_/Y input24/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0850_/X sky130_fd_sc_hd__mux2_2
XFILLER_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0781_ _1078_/Q _0777_/X input92/X _0778_/X vssd1 vssd1 vccd1 vccd1 _1078_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0755__A2 _0749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 addr_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0979_ _0978_/X _0979_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0979_/X sky130_fd_sc_hd__mux2_1
Xoutput363 _1037_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[50] sky130_fd_sc_hd__buf_2
Xoutput341 _1017_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[30] sky130_fd_sc_hd__buf_2
Xoutput352 _1027_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[40] sky130_fd_sc_hd__buf_2
Xoutput330 _1007_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[20] sky130_fd_sc_hd__buf_2
Xoutput385 _1057_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[70] sky130_fd_sc_hd__buf_2
Xoutput396 _1067_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[80] sky130_fd_sc_hd__buf_2
XFILLER_10_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput374 _1047_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[60] sky130_fd_sc_hd__buf_2
XFILLER_51_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input63_A data_to_core_mem[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0833_ _1114_/Q _0804_/A input97/X _0805_/A vssd1 vssd1 vccd1 vccd1 _1114_/D sky130_fd_sc_hd__a22o_1
X_0902_ _0902_/A0 _0902_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0902_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0764_ _0778_/A vssd1 vssd1 vccd1 vccd1 _0764_/X sky130_fd_sc_hd__clkbuf_2
X_0695_ _1019_/Q _0691_/X input73/X _0694_/X vssd1 vssd1 vccd1 vccd1 _1019_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0557__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0664__B2 _0659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0719__A2 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0655__B2 _0652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input215_A wr_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1101_ _1107_/CLK _1101_/D vssd1 vssd1 vccd1 vccd1 _1101_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0894__A1 _0894_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1032_ _1110_/CLK _1032_/D vssd1 vssd1 vccd1 vccd1 _1032_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0646__B2 _0645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput84 dout0_to_sram[1] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_4
X_0816_ _1101_/Q _0811_/X input82/X _0812_/X vssd1 vssd1 vccd1 vccd1 _1101_/D sky130_fd_sc_hd__a22o_1
Xinput95 dout0_to_sram[2] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_4
Xinput62 data_to_core_mem[29] vssd1 vssd1 vccd1 vccd1 _0633_/B sky130_fd_sc_hd__clkbuf_1
X_0747_ _1054_/Q _0740_/X input98/X _0743_/X vssd1 vssd1 vccd1 vccd1 _1054_/D sky130_fd_sc_hd__a22o_1
Xinput73 dout0_to_sram[0] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_2
Xinput40 addr_to_core_mem[9] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
Xinput51 data_to_core_mem[19] vssd1 vssd1 vccd1 vccd1 _0613_/B sky130_fd_sc_hd__clkbuf_1
X_0678_ _1011_/Q _0672_/X input89/X _0673_/X vssd1 vssd1 vccd1 vccd1 _1011_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0986__S _0986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0885__A1 _0884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0896__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input165_A wr_data[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0876__A1 _0876_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A addr_to_core_mem[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0800__A1 _1089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0601_ _0857_/S _0601_/B vssd1 vssd1 vccd1 vccd1 _0602_/A sky130_fd_sc_hd__and2_1
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0532_ _0532_/A vssd1 vssd1 vccd1 vccd1 _0532_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1015_ _1106_/CLK _1015_/D vssd1 vssd1 vccd1 vccd1 _1015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0858__A1 _0858_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0794__B1 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput230 wr_data[93] vssd1 vssd1 vccd1 vccd1 _0974_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__0849__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0785__B1 input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0515_ _0513_/A _0511_/Y _0517_/A vssd1 vssd1 vccd1 vccd1 _0515_/X sky130_fd_sc_hd__o21a_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0776__B1 input89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input128_A wr_data[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input93_A dout0_to_sram[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0767__B1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0995_ _1116_/CLK _0995_/D vssd1 vssd1 vccd1 vccd1 _0995_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0758__B1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0930__A0 _0930_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0780_ _1077_/Q _0777_/X input91/X _0778_/X vssd1 vssd1 vccd1 vccd1 _1077_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput5 addr_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
XANTENNA__0912__A0 _0911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0978_ _0978_/A0 _0978_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0978_/X sky130_fd_sc_hd__mux2_1
Xoutput331 _1008_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[21] sky130_fd_sc_hd__buf_2
Xoutput386 _1058_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[71] sky130_fd_sc_hd__buf_2
Xoutput364 _1038_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[51] sky130_fd_sc_hd__buf_2
Xoutput375 _1048_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[61] sky130_fd_sc_hd__buf_2
Xoutput320 _1114_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[127] sky130_fd_sc_hd__buf_2
Xoutput342 _1018_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[31] sky130_fd_sc_hd__buf_2
Xoutput397 _1068_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[81] sky130_fd_sc_hd__buf_2
Xoutput353 _1028_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[41] sky130_fd_sc_hd__buf_2
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input195_A wr_data[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A data_to_core_mem[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0899__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0901_ _0596_/X _0900_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1132_/D sky130_fd_sc_hd__mux2_1
X_0832_ _1113_/Q _0804_/A input96/X _0805_/A vssd1 vssd1 vccd1 vccd1 _1113_/D sky130_fd_sc_hd__a22o_1
X_0763_ _0777_/A vssd1 vssd1 vccd1 vccd1 _0763_/X sky130_fd_sc_hd__clkbuf_2
X_0694_ _0708_/A vssd1 vssd1 vccd1 vccd1 _0694_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0664__A2 _0658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input110_A wr_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0655__A2 _0651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input208_A wr_data[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_clk clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 _1109_/CLK sky130_fd_sc_hd__clkbuf_2
X_1100_ _1100_/CLK _1100_/D vssd1 vssd1 vccd1 vccd1 _1100_/Q sky130_fd_sc_hd__dfxtp_1
X_1031_ _1110_/CLK _1031_/D vssd1 vssd1 vccd1 vccd1 _1031_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0646__A2 _0642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0815_ _1100_/Q _0811_/X input81/X _0812_/X vssd1 vssd1 vccd1 vccd1 _1100_/D sky130_fd_sc_hd__a22o_1
Xinput30 addr_to_core_mem[18] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
Xinput41 data_to_core_mem[0] vssd1 vssd1 vccd1 vccd1 _0566_/A sky130_fd_sc_hd__clkbuf_1
Xinput96 dout0_to_sram[30] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__buf_2
XANTENNA__1149__GATE_N _0834_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0746_ _1053_/Q _0740_/X input95/X _0743_/X vssd1 vssd1 vccd1 vccd1 _1053_/D sky130_fd_sc_hd__a22o_1
Xinput74 dout0_to_sram[10] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_4
Xinput85 dout0_to_sram[20] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__buf_4
Xinput63 data_to_core_mem[2] vssd1 vssd1 vccd1 vccd1 _0579_/B sky130_fd_sc_hd__clkbuf_1
Xinput52 data_to_core_mem[1] vssd1 vssd1 vccd1 vccd1 _0577_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0677_ _1010_/Q _0672_/X input88/X _0673_/X vssd1 vssd1 vccd1 vccd1 _1010_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input158_A wr_data[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A addr_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0600_ _0600_/A vssd1 vssd1 vccd1 vccd1 _0600_/X sky130_fd_sc_hd__clkbuf_2
X_0531_ input2/X vssd1 vssd1 vccd1 vccd1 _0536_/A sky130_fd_sc_hd__inv_2
XANTENNA_output377_A _1050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1150__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1014_ _1112_/CLK _1014_/D vssd1 vssd1 vccd1 vccd1 _1014_/Q sky130_fd_sc_hd__dfxtp_1
X_0729_ _0729_/A vssd1 vssd1 vccd1 vccd1 _0729_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0794__B2 _0791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput231 wr_data[94] vssd1 vssd1 vccd1 vccd1 _0978_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput220 wr_data[84] vssd1 vssd1 vccd1 vccd1 _0938_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0514_ _0522_/A _0522_/B _0522_/D vssd1 vssd1 vccd1 vccd1 _0517_/A sky130_fd_sc_hd__or3_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0581__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0776__B2 _0771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input86_A dout0_to_sram[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output242_A _0851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0994_ _1065_/CLK _0994_/D vssd1 vssd1 vccd1 vccd1 _0994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input140_A wr_data[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0685__B1 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 addr_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0676__B1 input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput310 _1105_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[118] sky130_fd_sc_hd__buf_2
Xoutput332 _1009_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[22] sky130_fd_sc_hd__buf_2
X_0977_ _0634_/X _0976_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1151_/D sky130_fd_sc_hd__mux2_1
Xoutput321 _0999_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[12] sky130_fd_sc_hd__buf_2
Xoutput343 _1019_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[32] sky130_fd_sc_hd__buf_2
Xoutput354 _1029_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[42] sky130_fd_sc_hd__buf_2
Xoutput365 _1039_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[52] sky130_fd_sc_hd__buf_2
Xoutput376 _1049_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[62] sky130_fd_sc_hd__buf_2
XFILLER_19_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput398 _1069_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[82] sky130_fd_sc_hd__buf_2
Xoutput387 _1059_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[72] sky130_fd_sc_hd__buf_2
XANTENNA__0667__B1 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input188_A wr_data[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input49_A data_to_core_mem[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0900_ _0899_/X _0900_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0900_/X sky130_fd_sc_hd__mux2_2
X_0693_ _0729_/A vssd1 vssd1 vccd1 vccd1 _0708_/A sky130_fd_sc_hd__buf_2
X_0762_ _1065_/Q _0756_/X input78/X _0757_/X vssd1 vssd1 vccd1 vccd1 _1065_/D sky130_fd_sc_hd__a22o_1
X_0831_ _1112_/Q _0825_/X input94/X _0826_/X vssd1 vssd1 vccd1 vccd1 _1112_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0830__B1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1145__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0649__B1 input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0821__B1 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input103_A dout0_to_sram[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1030_ _1110_/CLK _1030_/D vssd1 vssd1 vccd1 vccd1 _1030_/Q sky130_fd_sc_hd__dfxtp_1
Xinput20 addr_in[9] vssd1 vssd1 vccd1 vccd1 _0528_/A sky130_fd_sc_hd__buf_2
XANTENNA__0803__B1 _0803_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput31 addr_to_core_mem[19] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
X_0814_ _1099_/Q _0811_/X input80/X _0812_/X vssd1 vssd1 vccd1 vccd1 _1099_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput86 dout0_to_sram[21] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_4
Xinput75 dout0_to_sram[11] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_4
Xinput97 dout0_to_sram[31] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_4
Xinput64 data_to_core_mem[30] vssd1 vssd1 vccd1 vccd1 _0635_/B sky130_fd_sc_hd__clkbuf_1
Xinput42 data_to_core_mem[10] vssd1 vssd1 vccd1 vccd1 _0595_/B sky130_fd_sc_hd__clkbuf_1
X_0676_ _1009_/Q _0672_/X input87/X _0673_/X vssd1 vssd1 vccd1 vccd1 _1009_/D sky130_fd_sc_hd__a22o_1
X_0745_ _1052_/Q _0740_/X input84/X _0743_/X vssd1 vssd1 vccd1 vccd1 _1052_/D sky130_fd_sc_hd__a22o_1
Xinput53 data_to_core_mem[20] vssd1 vssd1 vccd1 vccd1 _0615_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__0568__B _0568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input220_A wr_data[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0530_ _0528_/A _0526_/Y _0532_/A vssd1 vssd1 vccd1 vccd1 _0530_/X sky130_fd_sc_hd__o21a_2
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1013_ _1112_/CLK _1013_/D vssd1 vssd1 vccd1 vccd1 _1013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0728_ _0728_/A vssd1 vssd1 vccd1 vccd1 _0728_/X sky130_fd_sc_hd__clkbuf_2
X_0659_ _0659_/A vssd1 vssd1 vccd1 vccd1 _0659_/X sky130_fd_sc_hd__buf_2
XANTENNA__0579__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_clk clkbuf_4_9_0_clk/A vssd1 vssd1 vccd1 vccd1 _1111_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__0794__A2 _0788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input170_A wr_data[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput221 wr_data[85] vssd1 vssd1 vccd1 vccd1 _0942_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput232 wr_data[95] vssd1 vssd1 vccd1 vccd1 _0982_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input31_A addr_to_core_mem[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput210 wr_data[75] vssd1 vssd1 vccd1 vccd1 _0902_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0513_ _0513_/A vssd1 vssd1 vccd1 vccd1 _0522_/B sky130_fd_sc_hd__inv_2
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0776__A2 _0770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input79_A dout0_to_sram[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0993_ _1111_/CLK _0993_/D vssd1 vssd1 vccd1 vccd1 _0993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input133_A wr_data[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0685__A1 _1016_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput7 addr_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0676__B2 _0673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0976_ _0975_/X _0976_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0976_/X sky130_fd_sc_hd__mux2_2
Xoutput344 _1020_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[33] sky130_fd_sc_hd__buf_2
Xoutput355 _1030_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[43] sky130_fd_sc_hd__buf_2
Xoutput377 _1050_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[63] sky130_fd_sc_hd__buf_2
Xoutput322 _1000_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__1141__GATE_N _0834_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput300 _1096_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[109] sky130_fd_sc_hd__buf_2
Xoutput333 _1010_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[23] sky130_fd_sc_hd__buf_2
Xoutput366 _1040_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[53] sky130_fd_sc_hd__buf_2
Xoutput311 _1106_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[119] sky130_fd_sc_hd__buf_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput399 _1070_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[83] sky130_fd_sc_hd__buf_2
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput388 _1060_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[73] sky130_fd_sc_hd__buf_2
XANTENNA__0587__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0667__B2 _0666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0830__B2 _0826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0830_ _1111_/Q _0825_/X input93/X _0826_/X vssd1 vssd1 vccd1 vccd1 _1111_/D sky130_fd_sc_hd__a22o_1
X_0692_ _0728_/A vssd1 vssd1 vccd1 vccd1 _0729_/A sky130_fd_sc_hd__inv_2
X_0761_ _1064_/Q _0756_/X input77/X _0757_/X vssd1 vssd1 vccd1 vccd1 _1064_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0649__B2 _0645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0821__A1 _1104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0821__B2 _0819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0959_ _0958_/X _0959_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0959_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input61_A data_to_core_mem[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 addr_to_core_mem[0] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput43 data_to_core_mem[11] vssd1 vssd1 vccd1 vccd1 _0597_/B sky130_fd_sc_hd__buf_2
Xinput54 data_to_core_mem[21] vssd1 vssd1 vccd1 vccd1 _0617_/B sky130_fd_sc_hd__clkbuf_1
Xinput10 addr_in[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_2
X_0813_ _1098_/Q _0811_/X input79/X _0812_/X vssd1 vssd1 vccd1 vccd1 _1098_/D sky130_fd_sc_hd__a22o_1
Xinput32 addr_to_core_mem[1] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput65 data_to_core_mem[31] vssd1 vssd1 vccd1 vccd1 _0637_/B sky130_fd_sc_hd__clkbuf_1
X_0744_ _1051_/Q _0740_/X input73/X _0743_/X vssd1 vssd1 vccd1 vccd1 _1051_/D sky130_fd_sc_hd__a22o_1
X_0675_ _1008_/Q _0672_/X input86/X _0673_/X vssd1 vssd1 vccd1 vccd1 _1008_/D sky130_fd_sc_hd__a22o_1
Xinput76 dout0_to_sram[12] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_4
Xinput87 dout0_to_sram[22] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_4
Xinput98 dout0_to_sram[3] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1089_ _1107_/CLK _1089_/D vssd1 vssd1 vccd1 vccd1 _1089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0730__B1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input213_A wr_data[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1012_ _1106_/CLK _1012_/D vssd1 vssd1 vccd1 vccd1 _1012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0727_ _1043_/Q _0721_/X input89/X _0722_/X vssd1 vssd1 vccd1 vccd1 _1043_/D sky130_fd_sc_hd__a22o_1
X_0589_ _0857_/S _0589_/B vssd1 vssd1 vccd1 vccd1 _0590_/A sky130_fd_sc_hd__and2_1
X_0658_ _0658_/A vssd1 vssd1 vccd1 vccd1 _0658_/X sky130_fd_sc_hd__buf_2
XANTENNA__0595__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0712__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0779__B1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input163_A wr_data[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput233 wr_data[96] vssd1 vssd1 vccd1 vccd1 _0858_/A0 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input24_A addr_to_core_mem[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput222 wr_data[86] vssd1 vssd1 vccd1 vccd1 _0946_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput211 wr_data[76] vssd1 vssd1 vccd1 vccd1 _0906_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0703__B1 _0800_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput200 wr_data[66] vssd1 vssd1 vccd1 vccd1 _0866_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0942__A0 _0942_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0512_ _0522_/A _0522_/D _0511_/Y vssd1 vssd1 vccd1 vccd1 _0512_/Y sky130_fd_sc_hd__a21oi_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1136__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0924__A0 _0923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0992_ _1120_/CLK _0992_/D vssd1 vssd1 vccd1 vccd1 _0992_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0902__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_clk clkbuf_4_7_0_clk/A vssd1 vssd1 vccd1 vccd1 _1107_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input126_A wr_data[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input91_A dout0_to_sram[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 addr_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0676__A2 _0672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0975_ _0974_/X _0975_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0975_/X sky130_fd_sc_hd__mux2_1
Xoutput367 _1041_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[54] sky130_fd_sc_hd__buf_2
Xoutput378 _1051_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[64] sky130_fd_sc_hd__buf_2
Xoutput356 _1031_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[44] sky130_fd_sc_hd__buf_2
Xoutput301 _0997_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[10] sky130_fd_sc_hd__buf_2
Xoutput323 _1001_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[14] sky130_fd_sc_hd__buf_2
Xoutput334 _1011_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[24] sky130_fd_sc_hd__buf_2
Xoutput389 _1061_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[74] sky130_fd_sc_hd__buf_2
Xoutput312 _0998_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[11] sky130_fd_sc_hd__buf_2
Xoutput345 _1021_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[34] sky130_fd_sc_hd__buf_2
XANTENNA__0667__A2 _0665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0760_ _1063_/Q _0756_/X input76/X _0757_/X vssd1 vssd1 vccd1 vccd1 _1063_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0830__A2 _0825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0691_ _0707_/A vssd1 vssd1 vccd1 vccd1 _0691_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0649__A2 _0642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0889_ _0590_/X _0888_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1129_/D sky130_fd_sc_hd__mux2_4
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0958_ _0958_/A0 _0958_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0958_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input193_A wr_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input54_A data_to_core_mem[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput11 addr_in[19] vssd1 vssd1 vccd1 vccd1 _0564_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 addr_to_core_mem[10] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
Xinput55 data_to_core_mem[22] vssd1 vssd1 vccd1 vccd1 _0619_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput66 data_to_core_mem[3] vssd1 vssd1 vccd1 vccd1 _0581_/B sky130_fd_sc_hd__clkbuf_1
Xinput33 addr_to_core_mem[2] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0910__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput44 data_to_core_mem[12] vssd1 vssd1 vccd1 vccd1 _0599_/B sky130_fd_sc_hd__clkbuf_1
X_0743_ _0757_/A vssd1 vssd1 vccd1 vccd1 _0743_/X sky130_fd_sc_hd__buf_2
X_0812_ _0826_/A vssd1 vssd1 vccd1 vccd1 _0812_/X sky130_fd_sc_hd__buf_2
Xinput88 dout0_to_sram[23] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__buf_4
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput77 dout0_to_sram[13] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_4
Xinput99 dout0_to_sram[4] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__buf_2
X_0674_ _1007_/Q _0672_/X input85/X _0673_/X vssd1 vssd1 vccd1 vccd1 _1007_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1088_ _1107_/CLK _1088_/D vssd1 vssd1 vccd1 vccd1 _1088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input206_A wr_data[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1011_ _1112_/CLK _1011_/D vssd1 vssd1 vccd1 vccd1 _1011_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0905__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0726_ _1042_/Q _0721_/X input88/X _0722_/X vssd1 vssd1 vccd1 vccd1 _1042_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0712__B2 _0708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0657_ _0996_/Q _0651_/X _0803_/B1 _0652_/X vssd1 vssd1 vccd1 vccd1 _0996_/D sky130_fd_sc_hd__a22o_1
Xrepeater420 _0834_/Y vssd1 vssd1 vccd1 vccd1 repeater420/X sky130_fd_sc_hd__buf_12
X_0588_ _0588_/A vssd1 vssd1 vccd1 vccd1 _0588_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0951__A1 _0951_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1132__GATE_N _0834_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input156_A wr_data[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput201 wr_data[67] vssd1 vssd1 vccd1 vccd1 _0870_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput223 wr_data[87] vssd1 vssd1 vccd1 vccd1 _0950_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input17_A addr_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput212 wr_data[77] vssd1 vssd1 vccd1 vccd1 _0910_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput234 wr_data[97] vssd1 vssd1 vccd1 vccd1 _0862_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0511_ _0522_/A _0522_/D vssd1 vssd1 vccd1 vccd1 _0511_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0709_ _1029_/Q _0707_/X input74/X _0708_/X vssd1 vssd1 vccd1 vccd1 _1029_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0933__A1 _0932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input9_A addr_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0697__B1 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0991_ _1065_/CLK _0991_/D vssd1 vssd1 vccd1 vccd1 _0991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input119_A wr_data[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input84_A dout0_to_sram[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 addr_in[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0833__B1 input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0974_ _0974_/A0 _0974_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0974_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0913__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput313 _1107_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[120] sky130_fd_sc_hd__buf_2
Xoutput335 _1012_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[25] sky130_fd_sc_hd__buf_2
Xoutput324 _1002_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[15] sky130_fd_sc_hd__buf_2
Xoutput368 _1042_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[55] sky130_fd_sc_hd__buf_2
Xoutput302 _1097_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[110] sky130_fd_sc_hd__buf_2
XFILLER_19_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput357 _1032_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[45] sky130_fd_sc_hd__buf_2
Xoutput346 _1022_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[35] sky130_fd_sc_hd__buf_2
Xoutput379 _1052_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[65] sky130_fd_sc_hd__buf_2
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0824__B1 input89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input236_A wr_data[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0815__B1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_6_0_clk clkbuf_4_7_0_clk/A vssd1 vssd1 vccd1 vccd1 _1113_/CLK sky130_fd_sc_hd__clkbuf_2
X_0690_ _0728_/A vssd1 vssd1 vccd1 vccd1 _0707_/A sky130_fd_sc_hd__buf_2
XFILLER_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0908__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0806__B1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0957_ _0624_/X _0956_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1146_/D sky130_fd_sc_hd__mux2_2
X_0888_ _0887_/X _0888_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0888_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input47_A data_to_core_mem[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input186_A wr_data[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1127__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput78 dout0_to_sram[14] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__buf_4
Xinput56 data_to_core_mem[23] vssd1 vssd1 vccd1 vccd1 _0621_/B sky130_fd_sc_hd__clkbuf_1
X_0742_ _0778_/A vssd1 vssd1 vccd1 vccd1 _0757_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0811_ _0825_/A vssd1 vssd1 vccd1 vccd1 _0811_/X sky130_fd_sc_hd__buf_2
X_0673_ _0680_/A vssd1 vssd1 vccd1 vccd1 _0673_/X sky130_fd_sc_hd__buf_2
Xinput12 addr_in[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
Xinput45 data_to_core_mem[13] vssd1 vssd1 vccd1 vccd1 _0601_/B sky130_fd_sc_hd__clkbuf_1
Xinput23 addr_to_core_mem[11] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
Xinput34 addr_to_core_mem[3] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_2
Xinput89 dout0_to_sram[24] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_4
Xinput67 data_to_core_mem[4] vssd1 vssd1 vccd1 vccd1 _0583_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1087_ _1100_/CLK _1087_/D vssd1 vssd1 vccd1 vccd1 _1087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input101_A dout0_to_sram[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output418_A _0986_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1010_ _1094_/CLK _1010_/D vssd1 vssd1 vccd1 vccd1 _1010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0921__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0725_ _1041_/Q _0721_/X input87/X _0722_/X vssd1 vssd1 vccd1 vccd1 _1041_/D sky130_fd_sc_hd__a22o_1
X_0656_ _0995_/Q _0651_/X _0802_/B1 _0652_/X vssd1 vssd1 vccd1 vccd1 _0995_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0712__A2 _0707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0587_ _0857_/S _0587_/B vssd1 vssd1 vccd1 vccd1 _0588_/A sky130_fd_sc_hd__and2_1
X_1139_ _1139_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1139_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_4_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput213 wr_data[78] vssd1 vssd1 vccd1 vccd1 _0914_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput224 wr_data[88] vssd1 vssd1 vccd1 vccd1 _0954_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input149_A wr_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput202 wr_data[68] vssd1 vssd1 vccd1 vccd1 _0874_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput235 wr_data[98] vssd1 vssd1 vccd1 vccd1 _0866_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0510_ _0510_/A vssd1 vssd1 vccd1 vccd1 _0522_/A sky130_fd_sc_hd__inv_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0916__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0708_ _0708_/A vssd1 vssd1 vccd1 vccd1 _0708_/X sky130_fd_sc_hd__buf_2
X_0639_ _0568_/C _0568_/B _0857_/S vssd1 vssd1 vccd1 vccd1 _1121_/D sky130_fd_sc_hd__a21oi_1
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0990_ _1075_/CLK _0990_/D vssd1 vssd1 vccd1 vccd1 _0990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0851__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input77_A dout0_to_sram[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput303 _1098_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[111] sky130_fd_sc_hd__buf_2
X_0973_ _0632_/X _0972_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1150_/D sky130_fd_sc_hd__mux2_1
Xoutput314 _1108_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[121] sky130_fd_sc_hd__buf_2
Xoutput325 _1003_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[16] sky130_fd_sc_hd__buf_2
Xoutput369 _1043_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[56] sky130_fd_sc_hd__buf_2
Xoutput358 _1033_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[46] sky130_fd_sc_hd__buf_2
Xoutput347 _1023_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[36] sky130_fd_sc_hd__buf_2
Xoutput336 _1013_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0824__A1 _1107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0824__B2 _0819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input131_A wr_data[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0760__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input229_A wr_data[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0815__B2 _0812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1123__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0751__B1 _0799_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0956_ _0955_/X _0956_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0956_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0806__B2 _0805_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0924__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0887_ _0886_/X _0887_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0887_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0733__B1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input179_A wr_data[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 addr_in[2] vssd1 vssd1 vccd1 vccd1 _0501_/A sky130_fd_sc_hd__clkbuf_1
X_0810_ _1097_/Q _0804_/X input78/X _0805_/X vssd1 vssd1 vccd1 vccd1 _1097_/D sky130_fd_sc_hd__a22o_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput79 dout0_to_sram[15] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_4
Xinput24 addr_to_core_mem[12] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
Xinput57 data_to_core_mem[24] vssd1 vssd1 vccd1 vccd1 _0623_/B sky130_fd_sc_hd__clkbuf_1
Xinput68 data_to_core_mem[5] vssd1 vssd1 vccd1 vccd1 _0585_/B sky130_fd_sc_hd__clkbuf_1
X_0741_ _0777_/A vssd1 vssd1 vccd1 vccd1 _0778_/A sky130_fd_sc_hd__inv_2
X_0672_ _0679_/A vssd1 vssd1 vccd1 vccd1 _0672_/X sky130_fd_sc_hd__buf_2
Xinput46 data_to_core_mem[14] vssd1 vssd1 vccd1 vccd1 _0603_/B sky130_fd_sc_hd__clkbuf_1
Xinput35 addr_to_core_mem[4] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0919__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0724__B1 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1086_ _1113_/CLK _1086_/D vssd1 vssd1 vccd1 vccd1 _1086_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0939_ _0938_/X _0939_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0939_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5_0_clk clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 _1091_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0954__A0 _0954_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0706__B1 _0803_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output313_A _1107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0586_ _0586_/A vssd1 vssd1 vccd1 vccd1 _0586_/X sky130_fd_sc_hd__clkbuf_2
X_0724_ _1040_/Q _0721_/X input86/X _0722_/X vssd1 vssd1 vccd1 vccd1 _1040_/D sky130_fd_sc_hd__a22o_1
X_0655_ _0994_/Q _0651_/X _0801_/B1 _0652_/X vssd1 vssd1 vccd1 vccd1 _0994_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1138_ _1138_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1138_/Q sky130_fd_sc_hd__dlxtn_1
X_1069_ _1112_/CLK _1069_/D vssd1 vssd1 vccd1 vccd1 _1069_/Q sky130_fd_sc_hd__dfxtp_1
Xinput214 wr_data[79] vssd1 vssd1 vccd1 vccd1 _0918_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput203 wr_data[69] vssd1 vssd1 vccd1 vccd1 _0878_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput236 wr_data[99] vssd1 vssd1 vccd1 vccd1 _0870_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput225 wr_data[89] vssd1 vssd1 vccd1 vccd1 _0958_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input211_A wr_data[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0927__A0 _0926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0932__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0707_ _0707_/A vssd1 vssd1 vccd1 vccd1 _0707_/X sky130_fd_sc_hd__buf_2
XFILLER_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0638_ _0638_/A vssd1 vssd1 vccd1 vccd1 _0638_/X sky130_fd_sc_hd__clkbuf_1
X_0569_ _0569_/A vssd1 vssd1 vccd1 vccd1 _0985_/S sky130_fd_sc_hd__buf_12
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0842__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0909__A0 _0600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input161_A wr_data[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input22_A addr_to_core_mem[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0927__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0601__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0530__A1 _0528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0972_ _0971_/X _0972_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0972_/X sky130_fd_sc_hd__mux2_1
Xoutput359 _1034_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[47] sky130_fd_sc_hd__buf_2
Xoutput326 _1004_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[17] sky130_fd_sc_hd__buf_2
Xoutput315 _1109_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[122] sky130_fd_sc_hd__buf_2
Xoutput337 _1014_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[27] sky130_fd_sc_hd__buf_2
Xoutput304 _1099_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[112] sky130_fd_sc_hd__buf_2
Xoutput348 _1024_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[37] sky130_fd_sc_hd__buf_2
XFILLER_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input124_A wr_data[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0815__A2 _0811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0751__B2 _0750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output343_A _1019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0806__A2 _0804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0886_ _0886_/A0 _0886_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0886_/X sky130_fd_sc_hd__mux2_1
X_0955_ _0954_/X _0955_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0955_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0940__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0850__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0733__A1 _1047_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 addr_in[3] vssd1 vssd1 vccd1 vccd1 _0505_/A sky130_fd_sc_hd__clkbuf_1
Xinput25 addr_to_core_mem[13] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output293_A _1089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0740_ _0756_/A vssd1 vssd1 vccd1 vccd1 _0740_/X sky130_fd_sc_hd__buf_2
XFILLER_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput36 addr_to_core_mem[5] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput47 data_to_core_mem[15] vssd1 vssd1 vccd1 vccd1 _0605_/B sky130_fd_sc_hd__clkbuf_1
X_0671_ _1006_/Q _0665_/X input83/X _0666_/X vssd1 vssd1 vccd1 vccd1 _1006_/D sky130_fd_sc_hd__a22o_1
Xinput58 data_to_core_mem[25] vssd1 vssd1 vccd1 vccd1 _0625_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__0972__A1 _0972_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput69 data_to_core_mem[6] vssd1 vssd1 vccd1 vccd1 _0587_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__0724__B2 _0722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1085_ _1107_/CLK _1085_/D vssd1 vssd1 vccd1 vccd1 _1085_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0935__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0963__A1 _0963_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0869_ _0580_/X _0868_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1124_/D sky130_fd_sc_hd__mux2_1
X_0938_ _0938_/A0 _0938_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0938_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0660__B1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0845__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input191_A wr_data[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input52_A data_to_core_mem[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0890__A0 _0890_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0723_ _1039_/Q _0721_/X input85/X _0722_/X vssd1 vssd1 vccd1 vccd1 _1039_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0585_ _0857_/S _0585_/B vssd1 vssd1 vccd1 vccd1 _0586_/A sky130_fd_sc_hd__and2_1
X_0654_ _0993_/Q _0651_/X _0800_/B1 _0652_/X vssd1 vssd1 vccd1 vccd1 _0993_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1137_ _1137_/D _0834_/Y vssd1 vssd1 vccd1 vccd1 _1137_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0881__A0 _0586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1068_ _1112_/CLK _1068_/D vssd1 vssd1 vccd1 vccd1 _1068_/Q sky130_fd_sc_hd__dfxtp_1
Xinput204 wr_data[6] vssd1 vssd1 vccd1 vccd1 _0884_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput215 wr_data[7] vssd1 vssd1 vccd1 vccd1 _0888_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput237 wr_data[9] vssd1 vssd1 vccd1 vccd1 _0896_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput226 wr_data[8] vssd1 vssd1 vccd1 vccd1 _0892_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input204_A wr_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0927__A1 _0927_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_clk clkbuf_4_5_0_clk/A vssd1 vssd1 vccd1 vccd1 _1114_/CLK sky130_fd_sc_hd__clkbuf_2
X_0706_ _1028_/Q _0700_/X _0803_/B1 _0701_/X vssd1 vssd1 vccd1 vccd1 _1028_/D sky130_fd_sc_hd__a22o_1
X_0637_ _0857_/S _0637_/B vssd1 vssd1 vccd1 vccd1 _0638_/A sky130_fd_sc_hd__and2_1
X_0568_ _0857_/S _0568_/B _0568_/C vssd1 vssd1 vccd1 vccd1 _0569_/A sky130_fd_sc_hd__and3b_1
X_0499_ _1119_/Q input12/X _1119_/Q input12/X vssd1 vssd1 vccd1 vccd1 _0499_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input154_A wr_data[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input15_A addr_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0943__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input7_A addr_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0853__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_4_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0827__B1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1135__D _1135_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ _0970_/X _0971_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0971_/X sky130_fd_sc_hd__mux2_1
Xoutput305 _1100_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[113] sky130_fd_sc_hd__buf_2
Xoutput327 _1005_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[18] sky130_fd_sc_hd__buf_2
Xoutput316 _1110_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[123] sky130_fd_sc_hd__buf_2
Xoutput338 _1015_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[28] sky130_fd_sc_hd__buf_2
Xoutput349 _1025_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[38] sky130_fd_sc_hd__buf_2
XANTENNA__0938__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0809__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0848__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input117_A wr_data[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input82_A dout0_to_sram[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0751__A2 _0749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0954_ _0954_/A0 _0954_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0954_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0885_ _0588_/X _0884_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1128_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input234_A wr_data[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0607__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput59 data_to_core_mem[26] vssd1 vssd1 vccd1 vccd1 _0627_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 addr_to_core_mem[6] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
X_0670_ _1005_/Q _0665_/X input82/X _0666_/X vssd1 vssd1 vccd1 vccd1 _1005_/D sky130_fd_sc_hd__a22o_1
Xinput15 addr_in[4] vssd1 vssd1 vccd1 vccd1 _0510_/A sky130_fd_sc_hd__buf_2
Xinput26 addr_to_core_mem[14] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
Xinput48 data_to_core_mem[16] vssd1 vssd1 vccd1 vccd1 _0607_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0724__A2 _0721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1153_ _1153_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1153_/Q sky130_fd_sc_hd__dlxtn_1
X_1084_ _1107_/CLK _1084_/D vssd1 vssd1 vccd1 vccd1 _1084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0951__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0660__B2 _0659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0799_ _1088_/Q _0797_/X _0799_/B1 _0798_/X vssd1 vssd1 vccd1 vccd1 _1088_/D sky130_fd_sc_hd__a22o_1
X_0868_ _0867_/X _0868_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0868_/X sky130_fd_sc_hd__mux2_1
X_0937_ _0614_/X _0936_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1141_/D sky130_fd_sc_hd__mux2_2
XFILLER_57_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0861__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input45_A data_to_core_mem[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input184_A wr_data[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0722_ _0729_/A vssd1 vssd1 vccd1 vccd1 _0722_/X sky130_fd_sc_hd__buf_2
X_0653_ _0992_/Q _0651_/X _0799_/B1 _0652_/X vssd1 vssd1 vccd1 vccd1 _0992_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0584_ _0584_/A vssd1 vssd1 vccd1 vccd1 _0584_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0946__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1067_ _1106_/CLK _1067_/D vssd1 vssd1 vccd1 vccd1 _1067_/Q sky130_fd_sc_hd__dfxtp_1
X_1136_ _1136_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1136_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0856__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput205 wr_data[70] vssd1 vssd1 vccd1 vccd1 _0882_/A1 sky130_fd_sc_hd__buf_2
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput227 wr_data[90] vssd1 vssd1 vccd1 vccd1 _0962_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput216 wr_data[80] vssd1 vssd1 vccd1 vccd1 _0922_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output249_A _0839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output416_A _1086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0863__A1 _0863_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0636_ _0636_/A vssd1 vssd1 vccd1 vccd1 _0636_/X sky130_fd_sc_hd__clkbuf_1
X_0705_ _1027_/Q _0700_/X _0802_/B1 _0701_/X vssd1 vssd1 vccd1 vccd1 _1027_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0567_ _0567_/A vssd1 vssd1 vccd1 vccd1 _0567_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0498_ _0575_/D _0497_/B _0497_/Y vssd1 vssd1 vccd1 vccd1 _0498_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1119_ _1120_/CLK _1119_/D vssd1 vssd1 vccd1 vccd1 _1119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input147_A wr_data[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0615__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0781__B1 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0533__B1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0619_ _0857_/S _0619_/B vssd1 vssd1 vccd1 vccd1 _0620_/A sky130_fd_sc_hd__and2_1
XFILLER_49_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0772__B1 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0827__B2 _0826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_clk clkbuf_4_3_0_clk/A vssd1 vssd1 vccd1 vccd1 _1106_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0970_ _0970_/A0 _0970_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0970_/X sky130_fd_sc_hd__mux2_1
Xoutput306 _1101_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[114] sky130_fd_sc_hd__buf_2
Xoutput328 _1006_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[19] sky130_fd_sc_hd__buf_2
Xoutput317 _1111_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[124] sky130_fd_sc_hd__buf_2
Xoutput339 _1016_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[29] sky130_fd_sc_hd__buf_2
XANTENNA__0754__B1 _0802_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0954__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0809__B2 _0805_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0745__B1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0864__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0736__B1 input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input75_A dout0_to_sram[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1146__D _1146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0884_ _0883_/X _0884_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0884_/X sky130_fd_sc_hd__mux2_1
X_0953_ _0622_/X _0952_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1145_/D sky130_fd_sc_hd__mux2_1
XANTENNA__0727__B1 input89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0949__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0859__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0718__B1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input227_A wr_data[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput27 addr_to_core_mem[15] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0623__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput16 addr_in[5] vssd1 vssd1 vccd1 vccd1 _0513_/A sky130_fd_sc_hd__buf_2
Xinput38 addr_to_core_mem[7] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
Xinput49 data_to_core_mem[17] vssd1 vssd1 vccd1 vccd1 _0609_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0709__B1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1083_ _1083_/CLK _1083_/D vssd1 vssd1 vccd1 vccd1 _1083_/Q sky130_fd_sc_hd__dfxtp_2
X_1152_ _1152_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1152_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0936_ _0935_/X _0936_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0936_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0660__A2 _0658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0798_ _0805_/A vssd1 vssd1 vccd1 vccd1 _0798_/X sky130_fd_sc_hd__clkbuf_2
X_0867_ _0866_/X _0867_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0867_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0708__A _0708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input177_A wr_data[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input38_A addr_to_core_mem[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0721_ _0728_/A vssd1 vssd1 vccd1 vccd1 _0721_/X sky130_fd_sc_hd__buf_2
X_0652_ _0659_/A vssd1 vssd1 vccd1 vccd1 _0652_/X sky130_fd_sc_hd__clkbuf_4
X_0583_ _0857_/S _0583_/B vssd1 vssd1 vccd1 vccd1 _0584_/A sky130_fd_sc_hd__and2_1
XFILLER_6_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0962__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0528__A _0528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1135_ _1135_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1135_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1066_ _1106_/CLK _1066_/D vssd1 vssd1 vccd1 vccd1 _1066_/Q sky130_fd_sc_hd__dfxtp_1
X_0919_ _0918_/X _0919_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0919_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput206 wr_data[71] vssd1 vssd1 vccd1 vccd1 _0886_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput217 wr_data[81] vssd1 vssd1 vccd1 vccd1 _0926_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput228 wr_data[91] vssd1 vssd1 vccd1 vccd1 _0966_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0872__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output409_A _1079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0566_ _0566_/A _0857_/S vssd1 vssd1 vccd1 vccd1 _0567_/A sky130_fd_sc_hd__and2_1
X_0635_ _0857_/S _0635_/B vssd1 vssd1 vccd1 vccd1 _0636_/A sky130_fd_sc_hd__and2_1
X_0704_ _1026_/Q _0700_/X _0801_/B1 _0701_/X vssd1 vssd1 vccd1 vccd1 _1026_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0957__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0497_ _0575_/D _0497_/B vssd1 vssd1 vccd1 vccd1 _0497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1049_ _1100_/CLK _1049_/D vssd1 vssd1 vccd1 vccd1 _1049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1118_ _1120_/CLK _1118_/D vssd1 vssd1 vccd1 vccd1 _1118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0867__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1153__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0631__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0618_ _0618_/A vssd1 vssd1 vccd1 vccd1 _0618_/X sky130_fd_sc_hd__clkbuf_1
X_0549_ input7/X vssd1 vssd1 vccd1 vccd1 _0550_/B sky130_fd_sc_hd__inv_2
XANTENNA__0772__B2 _0771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0827__A2 _0825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0515__A1 _0513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input20_A addr_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput307 _1102_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[115] sky130_fd_sc_hd__buf_2
Xoutput329 _0988_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[1] sky130_fd_sc_hd__buf_2
Xoutput318 _1112_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[125] sky130_fd_sc_hd__buf_2
XANTENNA__0754__B2 _0750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0809__A2 _0804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0970__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0681__B1 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0984__A1 _0984_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0880__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0736__B2 _0708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0736__A1 _1050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input68_A data_to_core_mem[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0952_ _0951_/X _0952_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0952_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0883_ _0882_/X _0883_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0883_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0727__B2 _0722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0965__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0663__B1 input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_clk clkbuf_4_3_0_clk/A vssd1 vssd1 vccd1 vccd1 _1094_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__0718__B2 _0715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input122_A wr_data[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0875__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0654__B1 _0800_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 addr_in[6] vssd1 vssd1 vccd1 vccd1 _0516_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput28 addr_to_core_mem[16] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0709__B2 _0708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput39 addr_to_core_mem[8] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
X_1151_ _1151_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1151_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA_output341_A _1017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1082_ _1083_/CLK _1082_/D vssd1 vssd1 vccd1 vccd1 _1082_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0948__A1 _0948_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0935_ _0934_/X _0935_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0935_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0866_ _0866_/A0 _0866_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0866_/X sky130_fd_sc_hd__mux2_2
X_0797_ _0804_/A vssd1 vssd1 vccd1 vccd1 _0797_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0720_ _1038_/Q _0714_/X input83/X _0715_/X vssd1 vssd1 vccd1 vccd1 _1038_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0582_ _0582_/A vssd1 vssd1 vccd1 vccd1 _0582_/X sky130_fd_sc_hd__clkbuf_1
X_0651_ _0658_/A vssd1 vssd1 vccd1 vccd1 _0651_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1134_ _1134_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1134_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__1148__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1065_ _1065_/CLK _1065_/D vssd1 vssd1 vccd1 vccd1 _1065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0918_ _0918_/A0 _0918_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0918_/X sky130_fd_sc_hd__mux2_1
X_0849_ _0539_/X input23/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0849_/X sky130_fd_sc_hd__mux2_1
Xinput218 wr_data[82] vssd1 vssd1 vccd1 vccd1 _0930_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput207 wr_data[72] vssd1 vssd1 vccd1 vccd1 _0890_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput229 wr_data[92] vssd1 vssd1 vccd1 vccd1 _0970_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input50_A data_to_core_mem[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0629__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0703_ _1025_/Q _0700_/X _0800_/B1 _0701_/X vssd1 vssd1 vccd1 vccd1 _1025_/D sky130_fd_sc_hd__a22o_1
X_0565_ _0564_/A _0563_/A _0564_/Y _0561_/A vssd1 vssd1 vccd1 vccd1 _0565_/X sky130_fd_sc_hd__o22a_1
X_0634_ _0634_/A vssd1 vssd1 vccd1 vccd1 _0634_/X sky130_fd_sc_hd__clkbuf_1
X_0496_ input1/X vssd1 vssd1 vccd1 vccd1 _0497_/B sky130_fd_sc_hd__inv_2
XFILLER_53_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0973__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1117_ _1120_/CLK _1117_/D vssd1 vssd1 vccd1 vccd1 _1117_/Q sky130_fd_sc_hd__dfxtp_2
X_1048_ _1114_/CLK _1048_/D vssd1 vssd1 vccd1 vccd1 _1048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0883__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input202_A wr_data[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input98_A dout0_to_sram[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0772__A2 _0770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0617_ _0857_/S _0617_/B vssd1 vssd1 vccd1 vccd1 _0618_/A sky130_fd_sc_hd__and2_1
X_0548_ _0550_/A _0547_/A input6/X _0547_/Y vssd1 vssd1 vccd1 vccd1 _0548_/X sky130_fd_sc_hd__o22a_2
XANTENNA__0968__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0878__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input152_A wr_data[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A addr_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput308 _1103_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[116] sky130_fd_sc_hd__buf_2
Xoutput319 _1113_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[126] sky130_fd_sc_hd__buf_2
XANTENNA__0754__A2 _0749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A addr_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0736__A2 _0707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0637__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0882_ _0882_/A0 _0882_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0882_/X sky130_fd_sc_hd__mux2_1
X_0951_ _0950_/X _0951_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0951_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0727__A2 _0721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0981__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0663__B2 _0659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0718__A2 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input115_A wr_data[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput18 addr_in[7] vssd1 vssd1 vccd1 vccd1 _0519_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input80_A dout0_to_sram[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0654__B2 _0652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0891__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0709__A2 _0707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput29 addr_to_core_mem[17] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1150_ _1150_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1150_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1081_ _1083_/CLK _1081_/D vssd1 vssd1 vccd1 vccd1 _1081_/Q sky130_fd_sc_hd__dfxtp_1
X_0934_ _0934_/A0 _0934_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0934_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0865_ _0578_/X _0864_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1123_/D sky130_fd_sc_hd__mux2_2
X_0796_ _1087_/Q _0788_/X input99/X _0791_/X vssd1 vssd1 vccd1 vccd1 _1087_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1144__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0976__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0886__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input232_A wr_data[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0875__A1 _0875_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0581_ _0857_/S _0581_/B vssd1 vssd1 vccd1 vccd1 _0582_/A sky130_fd_sc_hd__and2_1
X_0650_ _0991_/Q _0642_/X input99/X _0645_/X vssd1 vssd1 vccd1 vccd1 _0991_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1064_ _1065_/CLK _1064_/D vssd1 vssd1 vccd1 vccd1 _1064_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_1_0_clk clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 _1110_/CLK sky130_fd_sc_hd__clkbuf_2
X_1133_ _1133_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1133_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0848_ _0533_/X input22/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0848_/X sky130_fd_sc_hd__mux2_4
X_0917_ _0604_/X _0916_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1136_/D sky130_fd_sc_hd__mux2_1
X_0779_ _1076_/Q _0777_/X input90/X _0778_/X vssd1 vssd1 vccd1 vccd1 _1076_/D sky130_fd_sc_hd__a22o_1
Xinput219 wr_data[83] vssd1 vssd1 vccd1 vccd1 _0934_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput208 wr_data[73] vssd1 vssd1 vccd1 vccd1 _0894_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0793__B1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input182_A wr_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A data_to_core_mem[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0633_ _0857_/S _0633_/B vssd1 vssd1 vccd1 vccd1 _0634_/A sky130_fd_sc_hd__and2_1
XANTENNA__0784__B1 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0702_ _1024_/Q _0700_/X _0799_/B1 _0701_/X vssd1 vssd1 vccd1 vccd1 _1024_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0564_ _0564_/A vssd1 vssd1 vccd1 vccd1 _0564_/Y sky130_fd_sc_hd__inv_2
X_0495_ _1117_/Q vssd1 vssd1 vccd1 vccd1 _0575_/D sky130_fd_sc_hd__clkinv_4
XANTENNA__0555__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1047_ _1109_/CLK _1047_/D vssd1 vssd1 vccd1 vccd1 _1047_/Q sky130_fd_sc_hd__dfxtp_2
X_1116_ _1116_/CLK _1119_/Q vssd1 vssd1 vccd1 vccd1 _1116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0775__B1 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0766__B1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output247_A _0856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0616_ _0616_/A vssd1 vssd1 vccd1 vccd1 _0616_/X sky130_fd_sc_hd__clkbuf_2
X_0547_ _0547_/A vssd1 vssd1 vccd1 vccd1 _0547_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0984__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0748__B1 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input145_A wr_data[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0894__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput309 _1104_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[117] sky130_fd_sc_hd__buf_2
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0978__A0 _0978_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0979__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0902__A0 _0902_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1139__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0889__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0881_ _0586_/X _0880_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1127_/D sky130_fd_sc_hd__mux2_1
X_0950_ _0950_/A0 _0950_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0950_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0663__A2 _0658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1140__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input108_A reset_mem_req vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0654__A2 _0651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 addr_in[8] vssd1 vssd1 vccd1 vccd1 _0525_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input73_A dout0_to_sram[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1080_ _1094_/CLK _1080_/D vssd1 vssd1 vccd1 vccd1 _1080_/Q sky130_fd_sc_hd__dfxtp_1
X_0795_ _1086_/Q _0788_/X input98/X _0791_/X vssd1 vssd1 vccd1 vccd1 _1086_/D sky130_fd_sc_hd__a22o_1
X_0933_ _0612_/X _0932_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1140_/D sky130_fd_sc_hd__mux2_1
X_0864_ _0863_/X _0864_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0864_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input225_A wr_data[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0580_ _0580_/A vssd1 vssd1 vccd1 vccd1 _0580_/X sky130_fd_sc_hd__clkbuf_1
X_1132_ _1132_/D _0834_/Y vssd1 vssd1 vccd1 vccd1 _1132_/Q sky130_fd_sc_hd__dlxtn_1
X_1063_ _1065_/CLK _1063_/D vssd1 vssd1 vccd1 vccd1 _1063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0916_ _0915_/X _0916_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0916_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0778_ _0778_/A vssd1 vssd1 vccd1 vccd1 _0778_/X sky130_fd_sc_hd__buf_2
X_0847_ _0530_/X input40/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0847_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput209 wr_data[74] vssd1 vssd1 vccd1 vccd1 _0898_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0793__B2 _0791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0545__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0897__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input175_A wr_data[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input36_A addr_to_core_mem[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0563_ _0563_/A _0563_/B vssd1 vssd1 vccd1 vccd1 _0563_/Y sky130_fd_sc_hd__nor2_1
X_0632_ _0632_/A vssd1 vssd1 vccd1 vccd1 _0632_/X sky130_fd_sc_hd__clkbuf_1
X_0701_ _0708_/A vssd1 vssd1 vccd1 vccd1 _0701_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0494_ _0494_/A vssd1 vssd1 vccd1 vccd1 _1117_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1046_ _1114_/CLK _1046_/D vssd1 vssd1 vccd1 vccd1 _1046_/Q sky130_fd_sc_hd__dfxtp_1
X_1115_ _1116_/CLK _1117_/Q vssd1 vssd1 vccd1 vccd1 _1115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0775__B2 _0771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0_clk clkbuf_4_1_0_clk/A vssd1 vssd1 vccd1 vccd1 _1112_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0546_ input6/X vssd1 vssd1 vccd1 vccd1 _0550_/A sky130_fd_sc_hd__inv_2
X_0615_ _0857_/S _0615_/B vssd1 vssd1 vccd1 vccd1 _0616_/A sky130_fd_sc_hd__and2_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1029_ _1109_/CLK _1029_/D vssd1 vssd1 vccd1 vccd1 _1029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0920__A1 _0920_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1135__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0684__B1 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input138_A wr_data[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0911__A1 _0911_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0675__B1 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clk/X sky130_fd_sc_hd__clkbuf_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0529_ _0537_/A _0537_/B _0537_/D vssd1 vssd1 vccd1 vccd1 _0532_/A sky130_fd_sc_hd__or3_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0657__B1 _0803_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0880_ _0879_/X _0880_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0880_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0648__B1 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0820__B1 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0639__B1 _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input66_A data_to_core_mem[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0932_ _0931_/X _0932_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0932_/X sky130_fd_sc_hd__mux2_2
X_0794_ _1085_/Q _0788_/X input95/X _0791_/X vssd1 vssd1 vccd1 vccd1 _1085_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0802__B1 _0802_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0863_ _0862_/X _0863_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0863_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input120_A wr_data[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input218_A wr_data[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1131_ _1131_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1131_/Q sky130_fd_sc_hd__dlxtn_1
X_1062_ _1116_/CLK _1062_/D vssd1 vssd1 vccd1 vccd1 _1062_/Q sky130_fd_sc_hd__dfxtp_1
X_0915_ _0914_/X _0915_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0915_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0777_ _0777_/A vssd1 vssd1 vccd1 vccd1 _0777_/X sky130_fd_sc_hd__buf_2
X_0846_ _0527_/Y input39/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0846_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0793__A2 _0788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput290 _0987_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[0] sky130_fd_sc_hd__buf_2
XANTENNA_input168_A wr_data[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input29_A addr_to_core_mem[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0700_ _0707_/A vssd1 vssd1 vccd1 vccd1 _0700_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0562_ input8/X input9/X _0554_/A input10/X vssd1 vssd1 vccd1 vccd1 _0563_/B sky130_fd_sc_hd__a31oi_1
X_0631_ _0857_/S _0631_/B vssd1 vssd1 vccd1 vccd1 _0632_/A sky130_fd_sc_hd__and2_1
X_1114_ _1114_/CLK _1114_/D vssd1 vssd1 vccd1 vccd1 _1114_/Q sky130_fd_sc_hd__dfxtp_1
X_0493_ _0492_/A _0986_/X vssd1 vssd1 vccd1 vccd1 _0494_/A sky130_fd_sc_hd__and2b_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1045_ _1114_/CLK _1045_/D vssd1 vssd1 vccd1 vccd1 _1045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0775__A2 _0770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0829_ _1110_/Q _0825_/X input92/X _0826_/X vssd1 vssd1 vccd1 vccd1 _1110_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1131__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0545_ input5/X _0541_/Y _0547_/A vssd1 vssd1 vccd1 vccd1 _0545_/X sky130_fd_sc_hd__o21a_1
X_0614_ _0614_/A vssd1 vssd1 vccd1 vccd1 _0614_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__0566__B _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1028_ _1094_/CLK _1028_/D vssd1 vssd1 vccd1 vccd1 _1028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input200_A wr_data[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input96_A dout0_to_sram[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0675__B2 _0673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0528_ _0528_/A vssd1 vssd1 vccd1 vccd1 _0537_/B sky130_fd_sc_hd__inv_2
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0577__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input150_A wr_data[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input11_A addr_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0487__A _0487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0657__B2 _0652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0648__B2 _0645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput190 wr_data[57] vssd1 vssd1 vccd1 vccd1 _0959_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0820__B2 _0819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input3_A addr_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input198_A wr_data[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input59_A data_to_core_mem[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_6_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0931_ _0930_/X _0931_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0931_/X sky130_fd_sc_hd__mux2_2
X_0862_ _0862_/A0 _0862_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0862_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0793_ _1084_/Q _0788_/X input84/X _0791_/X vssd1 vssd1 vccd1 vccd1 _1084_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input113_A wr_data[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0796__B1 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1126__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1130_ _1130_/D repeater420/X vssd1 vssd1 vccd1 vccd1 _1130_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__0720__B1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1061_ _1116_/CLK _1061_/D vssd1 vssd1 vccd1 vccd1 _1061_/Q sky130_fd_sc_hd__dfxtp_1
X_0914_ _0914_/A0 _0914_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0914_/X sky130_fd_sc_hd__mux2_1
X_0845_ _0524_/X input38/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0845_/X sky130_fd_sc_hd__mux2_2
X_0776_ _1075_/Q _0770_/X input89/X _0771_/X vssd1 vssd1 vccd1 vccd1 _1075_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0585__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0711__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput291 _1087_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[100] sky130_fd_sc_hd__buf_2
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input230_A wr_data[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput280 _1124_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[2] sky130_fd_sc_hd__buf_2
XANTENNA__0702__B1 _0799_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0769__B1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0561_ _0561_/A vssd1 vssd1 vccd1 vccd1 _0563_/A sky130_fd_sc_hd__inv_2
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0941__A0 _0616_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0630_ _0630_/A vssd1 vssd1 vccd1 vccd1 _0630_/X sky130_fd_sc_hd__clkbuf_1
X_0492_ _0492_/A _0492_/B vssd1 vssd1 vccd1 vccd1 _1118_/D sky130_fd_sc_hd__nor2_1
XFILLER_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1044_ _1083_/CLK _1044_/D vssd1 vssd1 vccd1 vccd1 _1044_/Q sky130_fd_sc_hd__dfxtp_1
X_1113_ _1113_/CLK _1113_/D vssd1 vssd1 vccd1 vccd1 _1113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0828_ _1109_/Q _0825_/X input91/X _0826_/X vssd1 vssd1 vccd1 vccd1 _1109_/D sky130_fd_sc_hd__a22o_1
X_0759_ _1062_/Q _0756_/X input75/X _0757_/X vssd1 vssd1 vccd1 vccd1 _1062_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0932__A0 _0931_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input41_A data_to_core_mem[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input180_A wr_data[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0613_ _0857_/S _0613_/B vssd1 vssd1 vccd1 vccd1 _0614_/A sky130_fd_sc_hd__and2_1
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0544_ _0551_/A _0551_/B _0551_/D vssd1 vssd1 vccd1 vccd1 _0547_/A sky130_fd_sc_hd__or3_2
XANTENNA__0914__A0 _0914_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1027_ _1094_/CLK _1027_/D vssd1 vssd1 vccd1 vccd1 _1027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input89_A dout0_to_sram[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0675__A2 _0672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0527_ _0537_/A _0537_/D _0526_/Y vssd1 vssd1 vccd1 vccd1 _0527_/Y sky130_fd_sc_hd__a21oi_4
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0593__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input143_A wr_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0487__B _0487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0657__A2 _0651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput180 wr_data[48] vssd1 vssd1 vccd1 vccd1 _0923_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0648__A2 _0642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput191 wr_data[58] vssd1 vssd1 vccd1 vccd1 _0963_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0639__A2 _0568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1122__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0861_ _0567_/X _0860_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1122_/D sky130_fd_sc_hd__mux2_1
X_0930_ _0930_/A0 _0930_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0930_/X sky130_fd_sc_hd__mux2_1
X_0792_ _1083_/Q _0788_/X input73/X _0791_/X vssd1 vssd1 vccd1 vccd1 _1083_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0900__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input106_A requested vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0796__B2 _0791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input71_A data_to_core_mem[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0720__B2 _0715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1060_ _1112_/CLK _1060_/D vssd1 vssd1 vccd1 vccd1 _1060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0691__A _0707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0844_ _0518_/X input37/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0844_/X sky130_fd_sc_hd__mux2_1
X_0775_ _1074_/Q _0770_/X input88/X _0771_/X vssd1 vssd1 vccd1 vccd1 _1074_/D sky130_fd_sc_hd__a22o_1
X_0913_ _0602_/X _0912_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1135_/D sky130_fd_sc_hd__mux2_2
XANTENNA__0711__B2 _0708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput270 _1142_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[20] sky130_fd_sc_hd__buf_2
Xclkbuf_3_5_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clk/X sky130_fd_sc_hd__clkbuf_2
Xoutput292 _1088_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[101] sky130_fd_sc_hd__buf_2
XANTENNA_input223_A wr_data[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput281 _1152_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[30] sky130_fd_sc_hd__buf_2
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0560_ _0560_/A _0560_/B _0560_/C input10/X vssd1 vssd1 vccd1 vccd1 _0561_/A sky130_fd_sc_hd__or4b_2
X_0491_ _1118_/Q _0485_/A _0575_/B _0571_/C vssd1 vssd1 vccd1 vccd1 _0492_/B sky130_fd_sc_hd__o22a_1
X_1043_ _1075_/CLK _1043_/D vssd1 vssd1 vccd1 vccd1 _1043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1112_ _1112_/CLK _1112_/D vssd1 vssd1 vccd1 vccd1 _1112_/Q sky130_fd_sc_hd__dfxtp_1
X_0758_ _1061_/Q _0756_/X input74/X _0757_/X vssd1 vssd1 vccd1 vccd1 _1061_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0827_ _1108_/Q _0825_/X input90/X _0826_/X vssd1 vssd1 vccd1 vccd1 _1108_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0596__A _0596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0689_ _0786_/A _1116_/Q vssd1 vssd1 vccd1 vccd1 _0728_/A sky130_fd_sc_hd__or2_2
XANTENNA__0696__B1 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input173_A wr_data[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0687__B1 input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A addr_to_core_mem[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0612_ _0612_/A vssd1 vssd1 vccd1 vccd1 _0612_/X sky130_fd_sc_hd__clkbuf_1
X_0543_ input5/X vssd1 vssd1 vccd1 vccd1 _0551_/B sky130_fd_sc_hd__inv_2
XFILLER_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0678__B1 input89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1026_ _1111_/CLK _1026_/D vssd1 vssd1 vccd1 vccd1 _1026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0669__B1 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output238_A _0838_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0832__B1 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0903__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0526_ _0537_/A _0537_/D vssd1 vssd1 vccd1 vccd1 _0526_/Y sky130_fd_sc_hd__nor2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1009_ _1091_/CLK _1009_/D vssd1 vssd1 vccd1 vccd1 _1009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0823__B1 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input136_A wr_data[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0814__B1 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output355_A _1030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput170 wr_data[39] vssd1 vssd1 vccd1 vccd1 _0887_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput181 wr_data[49] vssd1 vssd1 vccd1 vccd1 _0927_/A1 sky130_fd_sc_hd__buf_2
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput192 wr_data[59] vssd1 vssd1 vccd1 vccd1 _0967_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0694__A _0708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0509_ _0509_/A vssd1 vssd1 vccd1 vccd1 _0509_/X sky130_fd_sc_hd__clkbuf_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0860_ _0859_/X _0860_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0860_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0791_ _0805_/A vssd1 vssd1 vccd1 vccd1 _0791_/X sky130_fd_sc_hd__buf_2
XANTENNA_repeater420_A _0834_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0599__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0989_ _1113_/CLK _0989_/D vssd1 vssd1 vccd1 vccd1 _0989_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0796__A2 _0788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input64_A data_to_core_mem[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0720__A2 _0714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0912_ _0911_/X _0912_/A1 _0984_/S vssd1 vssd1 vccd1 vccd1 _0912_/X sky130_fd_sc_hd__mux2_1
X_0774_ _1073_/Q _0770_/X input87/X _0771_/X vssd1 vssd1 vccd1 vccd1 _1073_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0911__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0843_ _0515_/X input36/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0843_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0711__A2 _0707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput282 _1153_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[31] sky130_fd_sc_hd__buf_2
Xoutput271 _1143_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[21] sky130_fd_sc_hd__buf_2
Xoutput293 _1089_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[102] sky130_fd_sc_hd__buf_2
XFILLER_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput260 _1133_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[11] sky130_fd_sc_hd__buf_2
XFILLER_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input216_A wr_data[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0490_ _1118_/Q vssd1 vssd1 vccd1 vccd1 _0575_/B sky130_fd_sc_hd__inv_2
XFILLER_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1042_ _1075_/CLK _1042_/D vssd1 vssd1 vccd1 vccd1 _1042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0906__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1111_ _1111_/CLK _1111_/D vssd1 vssd1 vccd1 vccd1 _1111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0757_ _0757_/A vssd1 vssd1 vccd1 vccd1 _0757_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0688_ _1115_/Q vssd1 vssd1 vccd1 vccd1 _0786_/A sky130_fd_sc_hd__inv_2
X_0826_ _0826_/A vssd1 vssd1 vccd1 vccd1 _0826_/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _1075_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0696__A1 _1020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input166_A wr_data[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input27_A addr_to_core_mem[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0542_ _0551_/A _0551_/D _0541_/Y vssd1 vssd1 vccd1 vccd1 _0542_/Y sky130_fd_sc_hd__a21oi_1
X_0611_ _0857_/S _0611_/B vssd1 vssd1 vccd1 vccd1 _0612_/A sky130_fd_sc_hd__and2_1
XANTENNA__0678__B2 _0673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0850__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clk/A sky130_fd_sc_hd__clkbuf_2
X_1025_ _1111_/CLK _1025_/D vssd1 vssd1 vccd1 vccd1 _1025_/Q sky130_fd_sc_hd__dfxtp_1
X_0809_ _1096_/Q _0804_/X input77/X _0805_/X vssd1 vssd1 vccd1 vccd1 _1096_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0669__B2 _0666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0841__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0832__A1 _1113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0525_ _0525_/A vssd1 vssd1 vccd1 vccd1 _0537_/A sky130_fd_sc_hd__inv_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1008_ _1091_/CLK _1008_/D vssd1 vssd1 vccd1 vccd1 _1008_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0823__B2 _0819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input129_A wr_data[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input94_A dout0_to_sram[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0814__B2 _0812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output250_A _0840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput171 wr_data[3] vssd1 vssd1 vccd1 vccd1 _0872_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput182 wr_data[4] vssd1 vssd1 vccd1 vccd1 _0876_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput193 wr_data[5] vssd1 vssd1 vccd1 vccd1 _0880_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput160 wr_data[2] vssd1 vssd1 vccd1 vccd1 _0868_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA__0914__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0508_ _0506_/X _0522_/D vssd1 vssd1 vccd1 vccd1 _0509_/A sky130_fd_sc_hd__and2b_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0732__B1 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0799__B1 _0799_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0790_ _0826_/A vssd1 vssd1 vccd1 vccd1 _0805_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output298_A _1094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0723__B1 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0909__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0988_ _1065_/CLK _0988_/D vssd1 vssd1 vccd1 vccd1 _0988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input1_A addr_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input196_A wr_data[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input57_A data_to_core_mem[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0705__B1 _0802_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0911_ _0910_/X _0911_/A1 _0983_/S vssd1 vssd1 vccd1 vccd1 _0911_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0842_ _0512_/Y input35/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0842_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0773_ _1072_/Q _0770_/X input86/X _0771_/X vssd1 vssd1 vccd1 vccd1 _1072_/D sky130_fd_sc_hd__a22o_1
Xoutput294 _1090_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[103] sky130_fd_sc_hd__buf_2
Xoutput272 _1144_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[22] sky130_fd_sc_hd__buf_2
Xoutput283 _1125_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[3] sky130_fd_sc_hd__buf_2
Xoutput261 _1134_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[12] sky130_fd_sc_hd__buf_2
XANTENNA__0935__A0 _0934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput250 _0840_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[2] sky130_fd_sc_hd__buf_2
XANTENNA_input111_A wr_data[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input209_A wr_data[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1110_ _1110_/CLK _1110_/D vssd1 vssd1 vccd1 vccd1 _1110_/Q sky130_fd_sc_hd__dfxtp_1
X_1041_ _1075_/CLK _1041_/D vssd1 vssd1 vccd1 vccd1 _1041_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0922__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0825_ _0825_/A vssd1 vssd1 vccd1 vccd1 _0825_/X sky130_fd_sc_hd__buf_2
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0687_ _1018_/Q _0658_/A input97/X _0659_/A vssd1 vssd1 vccd1 vccd1 _1018_/D sky130_fd_sc_hd__a22o_1
X_0756_ _0756_/A vssd1 vssd1 vccd1 vccd1 _0756_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__0917__A0 _0604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input159_A wr_data[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output378_A _1051_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0541_ _0551_/A _0551_/D vssd1 vssd1 vccd1 vccd1 _0541_/Y sky130_fd_sc_hd__nor2_1
X_0610_ _0610_/A vssd1 vssd1 vccd1 vccd1 _0610_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1024_ _1094_/CLK _1024_/D vssd1 vssd1 vccd1 vccd1 _1024_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0678__A2 _0672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0917__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0835__C1 _0487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0808_ _1095_/Q _0804_/X input76/X _0805_/X vssd1 vssd1 vccd1 vccd1 _1095_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0669__A2 _0665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0739_ _0777_/A vssd1 vssd1 vccd1 vccd1 _0756_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _1065_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0524_ _0524_/A vssd1 vssd1 vccd1 vccd1 _0524_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1007_ _1112_/CLK _1007_/D vssd1 vssd1 vccd1 vccd1 _1007_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0814__A2 _0811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input87_A dout0_to_sram[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput161 wr_data[30] vssd1 vssd1 vccd1 vccd1 _0980_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput183 wr_data[50] vssd1 vssd1 vccd1 vccd1 _0931_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput194 wr_data[60] vssd1 vssd1 vccd1 vccd1 _0971_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput172 wr_data[40] vssd1 vssd1 vccd1 vccd1 _0891_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput150 wr_data[20] vssd1 vssd1 vccd1 vccd1 _0940_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_31_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0930__S _0982_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0507_ _0507_/A _0507_/B _0507_/C vssd1 vssd1 vccd1 vccd1 _0522_/D sky130_fd_sc_hd__or3_2
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0840__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input141_A wr_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output360_A _1035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0723__B2 _0722_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0925__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0987_ _1113_/CLK _0987_/D vssd1 vssd1 vccd1 vccd1 _0987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0962__A1 _0962_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput410 _1080_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[93] sky130_fd_sc_hd__buf_2
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0650__B1 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input189_A wr_data[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0910_ _0910_/A0 _0910_/A1 _0982_/S vssd1 vssd1 vccd1 vccd1 _0910_/X sky130_fd_sc_hd__mux2_1
X_0772_ _1071_/Q _0770_/X input85/X _0771_/X vssd1 vssd1 vccd1 vccd1 _1071_/D sky130_fd_sc_hd__a22o_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0841_ _0509_/X input34/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0841_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0944__A1 _0944_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0935__A1 _0935_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput273 _1145_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[23] sky130_fd_sc_hd__buf_2
Xoutput295 _1091_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[104] sky130_fd_sc_hd__buf_2
XFILLER_47_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput240 _0849_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[11] sky130_fd_sc_hd__buf_2
Xoutput251 _0841_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[3] sky130_fd_sc_hd__buf_2
Xoutput262 _1135_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[13] sky130_fd_sc_hd__buf_2
XANTENNA__0699__B1 input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput284 _1126_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[4] sky130_fd_sc_hd__buf_2
XANTENNA_input104_A dout0_to_sram[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1040_ _1065_/CLK _1040_/D vssd1 vssd1 vccd1 vccd1 _1040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0824_ _1107_/Q _0818_/X input89/X _0819_/X vssd1 vssd1 vccd1 vccd1 _1107_/D sky130_fd_sc_hd__a22o_1
XANTENNA__0917__A1 _0916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0755_ _1060_/Q _0749_/X _0803_/B1 _0750_/X vssd1 vssd1 vccd1 vccd1 _1060_/D sky130_fd_sc_hd__a22o_1
X_0686_ _1017_/Q _0658_/A input96/X _0659_/A vssd1 vssd1 vccd1 vccd1 _1017_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input221_A wr_data[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1130__D _1130_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0540_ input4/X vssd1 vssd1 vccd1 vccd1 _0551_/A sky130_fd_sc_hd__inv_2
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1023_ _1120_/CLK _1023_/D vssd1 vssd1 vccd1 vccd1 _1023_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__0835__B1 _0487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0933__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0738_ _1115_/Q _0786_/B vssd1 vssd1 vccd1 vccd1 _0777_/A sky130_fd_sc_hd__or2_2
X_0807_ _1094_/Q _0804_/X input75/X _0805_/X vssd1 vssd1 vccd1 vccd1 _1094_/D sky130_fd_sc_hd__a22o_1
X_0669_ _1004_/Q _0665_/X input81/X _0666_/X vssd1 vssd1 vccd1 vccd1 _1004_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0843__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input171_A wr_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input32_A addr_to_core_mem[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1152__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0817__B1 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0523_ _0520_/X _0537_/D vssd1 vssd1 vccd1 vccd1 _0524_/A sky130_fd_sc_hd__and2b_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0928__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1006_ _1091_/CLK _1006_/D vssd1 vssd1 vccd1 vccd1 _1006_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0808__B1 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0838__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput162 wr_data[31] vssd1 vssd1 vccd1 vccd1 _0984_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput151 wr_data[21] vssd1 vssd1 vccd1 vccd1 _0944_/A1 sky130_fd_sc_hd__buf_2
Xinput140 wr_data[127] vssd1 vssd1 vccd1 vccd1 _0982_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput173 wr_data[41] vssd1 vssd1 vccd1 vccd1 _0895_/A1 sky130_fd_sc_hd__buf_2
Xinput195 wr_data[61] vssd1 vssd1 vccd1 vccd1 _0975_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput184 wr_data[51] vssd1 vssd1 vccd1 vccd1 _0935_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0506_ _0507_/A _0507_/C _0507_/B vssd1 vssd1 vccd1 vccd1 _0506_/X sky130_fd_sc_hd__o21a_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _1100_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input134_A wr_data[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0723__A2 _0721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput400 _1071_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[84] sky130_fd_sc_hd__buf_2
Xoutput411 _1081_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[94] sky130_fd_sc_hd__buf_2
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0986_ _0575_/D _0568_/C _0986_/S vssd1 vssd1 vccd1 vccd1 _0986_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0941__S _0985_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0851__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0650__B2 _0645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0771_ _0778_/A vssd1 vssd1 vccd1 vccd1 _0771_/X sky130_fd_sc_hd__buf_2
X_0840_ _0504_/X input33/X _0857_/S vssd1 vssd1 vccd1 vccd1 _0840_/X sky130_fd_sc_hd__mux2_4
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__0936__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0880__A1 _0880_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0969_ _0630_/X _0968_/X _0985_/S vssd1 vssd1 vccd1 vccd1 _1149_/D sky130_fd_sc_hd__mux2_1
Xoutput252 _0842_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[4] sky130_fd_sc_hd__buf_2
Xoutput241 _0850_/X vssd1 vssd1 vccd1 vccd1 addr0_to_sram[12] sky130_fd_sc_hd__buf_2
Xoutput296 _1092_/Q vssd1 vssd1 vccd1 vccd1 rd_data_out[105] sky130_fd_sc_hd__buf_2
Xoutput285 _1127_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[5] sky130_fd_sc_hd__buf_2
Xoutput274 _1146_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[24] sky130_fd_sc_hd__buf_2
Xoutput263 _1136_/Q vssd1 vssd1 vccd1 vccd1 din0_to_sram[14] sky130_fd_sc_hd__buf_2
XANTENNA__0700__A _0707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0871__A1 _0871_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0846__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input62_A data_to_core_mem[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0754_ _1059_/Q _0749_/X _0802_/B1 _0750_/X vssd1 vssd1 vccd1 vccd1 _1059_/D sky130_fd_sc_hd__a22o_1
X_0685_ _1016_/Q _0679_/X input94/X _0680_/X vssd1 vssd1 vccd1 vccd1 _1016_/D sky130_fd_sc_hd__a22o_1
X_0823_ _1106_/Q _0818_/X input88/X _0819_/X vssd1 vssd1 vccd1 vccd1 _1106_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1147__GATE_N repeater420/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1099_ _1106_/CLK _1099_/D vssd1 vssd1 vccd1 vccd1 _1099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input214_A wr_data[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0605__A _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0780__B1 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1022_ _1120_/CLK _1022_/D vssd1 vssd1 vccd1 vccd1 _1022_/Q sky130_fd_sc_hd__dfxtp_1
X_0668_ _1003_/Q _0665_/X input80/X _0666_/X vssd1 vssd1 vccd1 vccd1 _1003_/D sky130_fd_sc_hd__a22o_1
X_0737_ _1116_/Q vssd1 vssd1 vccd1 vccd1 _0786_/B sky130_fd_sc_hd__inv_2
X_0806_ _1093_/Q _0804_/X input74/X _0805_/X vssd1 vssd1 vccd1 vccd1 _1093_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0599_ _0857_/S _0599_/B vssd1 vssd1 vccd1 vccd1 _0600_/A sky130_fd_sc_hd__and2_1
XFILLER_37_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0762__B1 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input164_A wr_data[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1141__D _1141_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_A addr_to_core_mem[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0817__B2 _0812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0522_ _0522_/A _0522_/B _0522_/C _0522_/D vssd1 vssd1 vccd1 vccd1 _0537_/D sky130_fd_sc_hd__or4_4
XANTENNA__0753__B1 _0801_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0944__S _0984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1005_ _1091_/CLK _1005_/D vssd1 vssd1 vccd1 vccd1 _1005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0808__B2 _0805_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0744__B1 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0854__S _0857_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0983__A0 _0982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0735__B1 input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput130 wr_data[118] vssd1 vssd1 vccd1 vccd1 _0946_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput141 wr_data[12] vssd1 vssd1 vccd1 vccd1 _0908_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput174 wr_data[42] vssd1 vssd1 vccd1 vccd1 _0899_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput152 wr_data[22] vssd1 vssd1 vccd1 vccd1 _0948_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput185 wr_data[52] vssd1 vssd1 vccd1 vccd1 _0939_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput163 wr_data[32] vssd1 vssd1 vccd1 vccd1 _0859_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput196 wr_data[62] vssd1 vssd1 vccd1 vccd1 _0979_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0505_ _0505_/A vssd1 vssd1 vccd1 vccd1 _0507_/B sky130_fd_sc_hd__inv_2
XANTENNA__0726__B1 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0939__S _0983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

