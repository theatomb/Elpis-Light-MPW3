VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO datapath
  CLASS BLOCK ;
  FOREIGN datapath ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 796.000 394.130 800.000 ;
    END
  END clk
  PIN current_address_rm2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 408.040 800.000 408.640 ;
    END
  END current_address_rm2[0]
  PIN current_address_rm2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 796.000 21.530 800.000 ;
    END
  END current_address_rm2[10]
  PIN current_address_rm2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END current_address_rm2[11]
  PIN current_address_rm2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END current_address_rm2[12]
  PIN current_address_rm2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 796.000 71.210 800.000 ;
    END
  END current_address_rm2[13]
  PIN current_address_rm2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 796.000 178.850 800.000 ;
    END
  END current_address_rm2[14]
  PIN current_address_rm2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END current_address_rm2[15]
  PIN current_address_rm2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 796.000 518.330 800.000 ;
    END
  END current_address_rm2[16]
  PIN current_address_rm2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 796.000 29.810 800.000 ;
    END
  END current_address_rm2[17]
  PIN current_address_rm2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END current_address_rm2[18]
  PIN current_address_rm2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 796.000 336.170 800.000 ;
    END
  END current_address_rm2[19]
  PIN current_address_rm2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 796.000 783.290 800.000 ;
    END
  END current_address_rm2[1]
  PIN current_address_rm2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END current_address_rm2[20]
  PIN current_address_rm2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 796.000 253.370 800.000 ;
    END
  END current_address_rm2[21]
  PIN current_address_rm2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 796.000 129.170 800.000 ;
    END
  END current_address_rm2[22]
  PIN current_address_rm2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 796.000 377.570 800.000 ;
    END
  END current_address_rm2[23]
  PIN current_address_rm2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 126.520 800.000 127.120 ;
    END
  END current_address_rm2[24]
  PIN current_address_rm2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END current_address_rm2[25]
  PIN current_address_rm2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END current_address_rm2[26]
  PIN current_address_rm2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 796.000 766.730 800.000 ;
    END
  END current_address_rm2[27]
  PIN current_address_rm2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.250 796.000 642.530 800.000 ;
    END
  END current_address_rm2[28]
  PIN current_address_rm2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 796.000 269.930 800.000 ;
    END
  END current_address_rm2[29]
  PIN current_address_rm2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 187.720 800.000 188.320 ;
    END
  END current_address_rm2[2]
  PIN current_address_rm2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 796.000 311.330 800.000 ;
    END
  END current_address_rm2[30]
  PIN current_address_rm2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 310.120 800.000 310.720 ;
    END
  END current_address_rm2[31]
  PIN current_address_rm2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 151.000 800.000 151.600 ;
    END
  END current_address_rm2[3]
  PIN current_address_rm2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END current_address_rm2[4]
  PIN current_address_rm2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 518.200 800.000 518.800 ;
    END
  END current_address_rm2[5]
  PIN current_address_rm2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END current_address_rm2[6]
  PIN current_address_rm2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 469.240 800.000 469.840 ;
    END
  END current_address_rm2[7]
  PIN current_address_rm2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END current_address_rm2[8]
  PIN current_address_rm2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END current_address_rm2[9]
  PIN dcache_re
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END dcache_re
  PIN exception_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END exception_type[0]
  PIN exception_type[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 796.000 410.690 800.000 ;
    END
  END exception_type[10]
  PIN exception_type[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 796.000 725.330 800.000 ;
    END
  END exception_type[11]
  PIN exception_type[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 175.480 800.000 176.080 ;
    END
  END exception_type[12]
  PIN exception_type[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END exception_type[13]
  PIN exception_type[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END exception_type[14]
  PIN exception_type[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 689.560 800.000 690.160 ;
    END
  END exception_type[15]
  PIN exception_type[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END exception_type[16]
  PIN exception_type[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 603.880 800.000 604.480 ;
    END
  END exception_type[17]
  PIN exception_type[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 616.120 800.000 616.720 ;
    END
  END exception_type[18]
  PIN exception_type[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 796.000 452.090 800.000 ;
    END
  END exception_type[19]
  PIN exception_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END exception_type[1]
  PIN exception_type[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 322.360 800.000 322.960 ;
    END
  END exception_type[20]
  PIN exception_type[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END exception_type[21]
  PIN exception_type[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 796.000 402.410 800.000 ;
    END
  END exception_type[22]
  PIN exception_type[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.650 796.000 683.930 800.000 ;
    END
  END exception_type[23]
  PIN exception_type[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END exception_type[24]
  PIN exception_type[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END exception_type[25]
  PIN exception_type[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 444.760 800.000 445.360 ;
    END
  END exception_type[26]
  PIN exception_type[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END exception_type[27]
  PIN exception_type[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 796.000 427.250 800.000 ;
    END
  END exception_type[28]
  PIN exception_type[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 763.000 800.000 763.600 ;
    END
  END exception_type[29]
  PIN exception_type[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 796.000 236.810 800.000 ;
    END
  END exception_type[2]
  PIN exception_type[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END exception_type[30]
  PIN exception_type[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END exception_type[31]
  PIN exception_type[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 796.000 286.490 800.000 ;
    END
  END exception_type[3]
  PIN exception_type[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 796.000 319.610 800.000 ;
    END
  END exception_type[4]
  PIN exception_type[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END exception_type[5]
  PIN exception_type[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 701.800 800.000 702.400 ;
    END
  END exception_type[6]
  PIN exception_type[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END exception_type[7]
  PIN exception_type[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 457.000 800.000 457.600 ;
    END
  END exception_type[8]
  PIN exception_type[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END exception_type[9]
  PIN hit_dcache
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END hit_dcache
  PIN hit_dtlb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END hit_dtlb
  PIN hit_icache
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END hit_icache
  PIN hit_itlb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END hit_itlb
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 796.000 54.650 800.000 ;
    END
  END is_print_done
  PIN is_read_interactive_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END is_read_interactive_enabled
  PIN is_tlbwrite
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 796.000 659.090 800.000 ;
    END
  END is_tlbwrite
  PIN mem_addr_f[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 796.000 584.570 800.000 ;
    END
  END mem_addr_f[0]
  PIN mem_addr_f[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 796.000 211.970 800.000 ;
    END
  END mem_addr_f[10]
  PIN mem_addr_f[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 796.000 38.090 800.000 ;
    END
  END mem_addr_f[11]
  PIN mem_addr_f[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END mem_addr_f[12]
  PIN mem_addr_f[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 224.440 800.000 225.040 ;
    END
  END mem_addr_f[13]
  PIN mem_addr_f[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 65.320 800.000 65.920 ;
    END
  END mem_addr_f[14]
  PIN mem_addr_f[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 796.000 700.490 800.000 ;
    END
  END mem_addr_f[15]
  PIN mem_addr_f[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 0.000 795.250 4.000 ;
    END
  END mem_addr_f[16]
  PIN mem_addr_f[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END mem_addr_f[17]
  PIN mem_addr_f[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 0.000 778.690 4.000 ;
    END
  END mem_addr_f[18]
  PIN mem_addr_f[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 796.000 534.890 800.000 ;
    END
  END mem_addr_f[19]
  PIN mem_addr_f[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 796.000 559.730 800.000 ;
    END
  END mem_addr_f[1]
  PIN mem_addr_f[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END mem_addr_f[20]
  PIN mem_addr_f[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 796.000 62.930 800.000 ;
    END
  END mem_addr_f[21]
  PIN mem_addr_f[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 796.000 617.690 800.000 ;
    END
  END mem_addr_f[22]
  PIN mem_addr_f[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END mem_addr_f[23]
  PIN mem_addr_f[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 796.000 791.570 800.000 ;
    END
  END mem_addr_f[24]
  PIN mem_addr_f[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 796.000 493.490 800.000 ;
    END
  END mem_addr_f[25]
  PIN mem_addr_f[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END mem_addr_f[26]
  PIN mem_addr_f[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END mem_addr_f[27]
  PIN mem_addr_f[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 796.000 327.890 800.000 ;
    END
  END mem_addr_f[28]
  PIN mem_addr_f[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 738.520 800.000 739.120 ;
    END
  END mem_addr_f[29]
  PIN mem_addr_f[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END mem_addr_f[2]
  PIN mem_addr_f[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END mem_addr_f[30]
  PIN mem_addr_f[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 796.000 460.370 800.000 ;
    END
  END mem_addr_f[31]
  PIN mem_addr_f[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 796.000 195.410 800.000 ;
    END
  END mem_addr_f[3]
  PIN mem_addr_f[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 796.000 187.130 800.000 ;
    END
  END mem_addr_f[4]
  PIN mem_addr_f[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END mem_addr_f[5]
  PIN mem_addr_f[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 212.200 800.000 212.800 ;
    END
  END mem_addr_f[6]
  PIN mem_addr_f[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END mem_addr_f[7]
  PIN mem_addr_f[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END mem_addr_f[8]
  PIN mem_addr_f[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END mem_addr_f[9]
  PIN mem_addr_m[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 796.000 162.290 800.000 ;
    END
  END mem_addr_m[0]
  PIN mem_addr_m[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END mem_addr_m[10]
  PIN mem_addr_m[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END mem_addr_m[11]
  PIN mem_addr_m[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END mem_addr_m[12]
  PIN mem_addr_m[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END mem_addr_m[13]
  PIN mem_addr_m[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 796.000 104.330 800.000 ;
    END
  END mem_addr_m[14]
  PIN mem_addr_m[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END mem_addr_m[15]
  PIN mem_addr_m[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END mem_addr_m[16]
  PIN mem_addr_m[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END mem_addr_m[17]
  PIN mem_addr_m[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 4.000 794.880 ;
    END
  END mem_addr_m[18]
  PIN mem_addr_m[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 796.000 543.170 800.000 ;
    END
  END mem_addr_m[19]
  PIN mem_addr_m[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END mem_addr_m[1]
  PIN mem_addr_m[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END mem_addr_m[20]
  PIN mem_addr_m[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 796.000 46.370 800.000 ;
    END
  END mem_addr_m[21]
  PIN mem_addr_m[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END mem_addr_m[22]
  PIN mem_addr_m[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END mem_addr_m[23]
  PIN mem_addr_m[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 493.720 800.000 494.320 ;
    END
  END mem_addr_m[24]
  PIN mem_addr_m[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 796.000 468.650 800.000 ;
    END
  END mem_addr_m[25]
  PIN mem_addr_m[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 371.320 800.000 371.920 ;
    END
  END mem_addr_m[26]
  PIN mem_addr_m[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END mem_addr_m[27]
  PIN mem_addr_m[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END mem_addr_m[28]
  PIN mem_addr_m[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END mem_addr_m[29]
  PIN mem_addr_m[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 796.000 4.970 800.000 ;
    END
  END mem_addr_m[2]
  PIN mem_addr_m[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 796.000 303.050 800.000 ;
    END
  END mem_addr_m[30]
  PIN mem_addr_m[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 579.400 800.000 580.000 ;
    END
  END mem_addr_m[31]
  PIN mem_addr_m[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END mem_addr_m[3]
  PIN mem_addr_m[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 796.000 385.850 800.000 ;
    END
  END mem_addr_m[4]
  PIN mem_addr_m[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END mem_addr_m[5]
  PIN mem_addr_m[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END mem_addr_m[6]
  PIN mem_addr_m[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END mem_addr_m[7]
  PIN mem_addr_m[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 89.800 800.000 90.400 ;
    END
  END mem_addr_m[8]
  PIN mem_addr_m[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END mem_addr_m[9]
  PIN mem_data_rd_f[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END mem_data_rd_f[0]
  PIN mem_data_rd_f[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 787.480 800.000 788.080 ;
    END
  END mem_data_rd_f[10]
  PIN mem_data_rd_f[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 114.280 800.000 114.880 ;
    END
  END mem_data_rd_f[11]
  PIN mem_data_rd_f[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 796.000 245.090 800.000 ;
    END
  END mem_data_rd_f[12]
  PIN mem_data_rd_f[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END mem_data_rd_f[13]
  PIN mem_data_rd_f[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.570 796.000 799.850 800.000 ;
    END
  END mem_data_rd_f[14]
  PIN mem_data_rd_f[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END mem_data_rd_f[15]
  PIN mem_data_rd_f[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 796.000 294.770 800.000 ;
    END
  END mem_data_rd_f[16]
  PIN mem_data_rd_f[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 0.000 563.410 4.000 ;
    END
  END mem_data_rd_f[17]
  PIN mem_data_rd_f[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END mem_data_rd_f[18]
  PIN mem_data_rd_f[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 420.280 800.000 420.880 ;
    END
  END mem_data_rd_f[19]
  PIN mem_data_rd_f[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END mem_data_rd_f[1]
  PIN mem_data_rd_f[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END mem_data_rd_f[20]
  PIN mem_data_rd_f[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END mem_data_rd_f[21]
  PIN mem_data_rd_f[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 163.240 800.000 163.840 ;
    END
  END mem_data_rd_f[22]
  PIN mem_data_rd_f[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END mem_data_rd_f[23]
  PIN mem_data_rd_f[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END mem_data_rd_f[24]
  PIN mem_data_rd_f[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 796.000 733.610 800.000 ;
    END
  END mem_data_rd_f[25]
  PIN mem_data_rd_f[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END mem_data_rd_f[26]
  PIN mem_data_rd_f[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END mem_data_rd_f[27]
  PIN mem_data_rd_f[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END mem_data_rd_f[28]
  PIN mem_data_rd_f[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END mem_data_rd_f[29]
  PIN mem_data_rd_f[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END mem_data_rd_f[2]
  PIN mem_data_rd_f[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 796.000 634.250 800.000 ;
    END
  END mem_data_rd_f[30]
  PIN mem_data_rd_f[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 40.840 800.000 41.440 ;
    END
  END mem_data_rd_f[31]
  PIN mem_data_rd_f[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END mem_data_rd_f[3]
  PIN mem_data_rd_f[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 542.680 800.000 543.280 ;
    END
  END mem_data_rd_f[4]
  PIN mem_data_rd_f[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 652.840 800.000 653.440 ;
    END
  END mem_data_rd_f[5]
  PIN mem_data_rd_f[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END mem_data_rd_f[6]
  PIN mem_data_rd_f[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 796.000 154.010 800.000 ;
    END
  END mem_data_rd_f[7]
  PIN mem_data_rd_f[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END mem_data_rd_f[8]
  PIN mem_data_rd_f[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 796.000 369.290 800.000 ;
    END
  END mem_data_rd_f[9]
  PIN mem_data_rd_m[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END mem_data_rd_m[0]
  PIN mem_data_rd_m[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END mem_data_rd_m[10]
  PIN mem_data_rd_m[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 432.520 800.000 433.120 ;
    END
  END mem_data_rd_m[11]
  PIN mem_data_rd_m[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 481.480 800.000 482.080 ;
    END
  END mem_data_rd_m[12]
  PIN mem_data_rd_m[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 359.080 800.000 359.680 ;
    END
  END mem_data_rd_m[13]
  PIN mem_data_rd_m[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 796.000 220.250 800.000 ;
    END
  END mem_data_rd_m[14]
  PIN mem_data_rd_m[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END mem_data_rd_m[15]
  PIN mem_data_rd_m[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END mem_data_rd_m[16]
  PIN mem_data_rd_m[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 591.640 800.000 592.240 ;
    END
  END mem_data_rd_m[17]
  PIN mem_data_rd_m[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 796.000 601.130 800.000 ;
    END
  END mem_data_rd_m[18]
  PIN mem_data_rd_m[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END mem_data_rd_m[19]
  PIN mem_data_rd_m[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 796.000 551.450 800.000 ;
    END
  END mem_data_rd_m[1]
  PIN mem_data_rd_m[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END mem_data_rd_m[20]
  PIN mem_data_rd_m[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 796.000 228.530 800.000 ;
    END
  END mem_data_rd_m[21]
  PIN mem_data_rd_m[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END mem_data_rd_m[22]
  PIN mem_data_rd_m[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END mem_data_rd_m[23]
  PIN mem_data_rd_m[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 796.000 625.970 800.000 ;
    END
  END mem_data_rd_m[24]
  PIN mem_data_rd_m[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END mem_data_rd_m[25]
  PIN mem_data_rd_m[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END mem_data_rd_m[26]
  PIN mem_data_rd_m[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END mem_data_rd_m[27]
  PIN mem_data_rd_m[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END mem_data_rd_m[28]
  PIN mem_data_rd_m[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END mem_data_rd_m[29]
  PIN mem_data_rd_m[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END mem_data_rd_m[2]
  PIN mem_data_rd_m[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END mem_data_rd_m[30]
  PIN mem_data_rd_m[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 102.040 800.000 102.640 ;
    END
  END mem_data_rd_m[31]
  PIN mem_data_rd_m[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 261.160 800.000 261.760 ;
    END
  END mem_data_rd_m[3]
  PIN mem_data_rd_m[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END mem_data_rd_m[4]
  PIN mem_data_rd_m[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END mem_data_rd_m[5]
  PIN mem_data_rd_m[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END mem_data_rd_m[6]
  PIN mem_data_rd_m[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 236.680 800.000 237.280 ;
    END
  END mem_data_rd_m[7]
  PIN mem_data_rd_m[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 796.000 775.010 800.000 ;
    END
  END mem_data_rd_m[8]
  PIN mem_data_rd_m[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 796.000 418.970 800.000 ;
    END
  END mem_data_rd_m[9]
  PIN mem_data_wr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END mem_data_wr[0]
  PIN mem_data_wr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 665.080 800.000 665.680 ;
    END
  END mem_data_wr[10]
  PIN mem_data_wr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END mem_data_wr[11]
  PIN mem_data_wr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END mem_data_wr[12]
  PIN mem_data_wr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END mem_data_wr[13]
  PIN mem_data_wr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END mem_data_wr[14]
  PIN mem_data_wr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END mem_data_wr[15]
  PIN mem_data_wr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 796.000 112.610 800.000 ;
    END
  END mem_data_wr[16]
  PIN mem_data_wr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 796.000 278.210 800.000 ;
    END
  END mem_data_wr[17]
  PIN mem_data_wr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 285.640 800.000 286.240 ;
    END
  END mem_data_wr[18]
  PIN mem_data_wr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END mem_data_wr[19]
  PIN mem_data_wr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END mem_data_wr[1]
  PIN mem_data_wr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 796.000 510.050 800.000 ;
    END
  END mem_data_wr[20]
  PIN mem_data_wr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 726.280 800.000 726.880 ;
    END
  END mem_data_wr[21]
  PIN mem_data_wr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 395.800 800.000 396.400 ;
    END
  END mem_data_wr[22]
  PIN mem_data_wr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 796.000 476.930 800.000 ;
    END
  END mem_data_wr[23]
  PIN mem_data_wr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 796.000 526.610 800.000 ;
    END
  END mem_data_wr[24]
  PIN mem_data_wr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END mem_data_wr[25]
  PIN mem_data_wr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 796.000 435.530 800.000 ;
    END
  END mem_data_wr[26]
  PIN mem_data_wr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 28.600 800.000 29.200 ;
    END
  END mem_data_wr[27]
  PIN mem_data_wr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 796.000 717.050 800.000 ;
    END
  END mem_data_wr[28]
  PIN mem_data_wr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 796.000 592.850 800.000 ;
    END
  END mem_data_wr[29]
  PIN mem_data_wr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END mem_data_wr[2]
  PIN mem_data_wr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END mem_data_wr[30]
  PIN mem_data_wr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 796.000 170.570 800.000 ;
    END
  END mem_data_wr[31]
  PIN mem_data_wr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 383.560 800.000 384.160 ;
    END
  END mem_data_wr[3]
  PIN mem_data_wr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END mem_data_wr[4]
  PIN mem_data_wr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END mem_data_wr[5]
  PIN mem_data_wr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 796.000 145.730 800.000 ;
    END
  END mem_data_wr[6]
  PIN mem_data_wr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 16.360 800.000 16.960 ;
    END
  END mem_data_wr[7]
  PIN mem_data_wr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END mem_data_wr[8]
  PIN mem_data_wr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 796.000 692.210 800.000 ;
    END
  END mem_data_wr[9]
  PIN mem_isbyte
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 714.040 800.000 714.640 ;
    END
  END mem_isbyte
  PIN mem_physical_tlb_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END mem_physical_tlb_addr_out[0]
  PIN mem_physical_tlb_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END mem_physical_tlb_addr_out[10]
  PIN mem_physical_tlb_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 0.000 762.130 4.000 ;
    END
  END mem_physical_tlb_addr_out[11]
  PIN mem_physical_tlb_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END mem_physical_tlb_addr_out[12]
  PIN mem_physical_tlb_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END mem_physical_tlb_addr_out[13]
  PIN mem_physical_tlb_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END mem_physical_tlb_addr_out[14]
  PIN mem_physical_tlb_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 796.000 485.210 800.000 ;
    END
  END mem_physical_tlb_addr_out[15]
  PIN mem_physical_tlb_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 273.400 800.000 274.000 ;
    END
  END mem_physical_tlb_addr_out[16]
  PIN mem_physical_tlb_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 628.360 800.000 628.960 ;
    END
  END mem_physical_tlb_addr_out[17]
  PIN mem_physical_tlb_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END mem_physical_tlb_addr_out[18]
  PIN mem_physical_tlb_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 796.000 758.450 800.000 ;
    END
  END mem_physical_tlb_addr_out[19]
  PIN mem_physical_tlb_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 138.760 800.000 139.360 ;
    END
  END mem_physical_tlb_addr_out[1]
  PIN mem_physical_tlb_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END mem_physical_tlb_addr_out[2]
  PIN mem_physical_tlb_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 796.000 741.890 800.000 ;
    END
  END mem_physical_tlb_addr_out[3]
  PIN mem_physical_tlb_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END mem_physical_tlb_addr_out[4]
  PIN mem_physical_tlb_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END mem_physical_tlb_addr_out[5]
  PIN mem_physical_tlb_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END mem_physical_tlb_addr_out[6]
  PIN mem_physical_tlb_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 0.000 629.650 4.000 ;
    END
  END mem_physical_tlb_addr_out[7]
  PIN mem_physical_tlb_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 4.120 800.000 4.720 ;
    END
  END mem_physical_tlb_addr_out[8]
  PIN mem_physical_tlb_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 796.000 443.810 800.000 ;
    END
  END mem_physical_tlb_addr_out[9]
  PIN mem_wrd
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 567.160 800.000 567.760 ;
    END
  END mem_wrd
  PIN print_hex_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 796.000 96.050 800.000 ;
    END
  END print_hex_enable
  PIN print_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 796.000 137.450 800.000 ;
    END
  END print_output[0]
  PIN print_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 796.000 120.890 800.000 ;
    END
  END print_output[10]
  PIN print_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END print_output[11]
  PIN print_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END print_output[12]
  PIN print_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 248.920 800.000 249.520 ;
    END
  END print_output[13]
  PIN print_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END print_output[14]
  PIN print_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 796.000 667.370 800.000 ;
    END
  END print_output[15]
  PIN print_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 775.240 800.000 775.840 ;
    END
  END print_output[16]
  PIN print_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 796.000 261.650 800.000 ;
    END
  END print_output[17]
  PIN print_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END print_output[18]
  PIN print_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END print_output[19]
  PIN print_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 750.760 800.000 751.360 ;
    END
  END print_output[1]
  PIN print_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END print_output[20]
  PIN print_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 505.960 800.000 506.560 ;
    END
  END print_output[21]
  PIN print_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END print_output[22]
  PIN print_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END print_output[23]
  PIN print_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 796.000 750.170 800.000 ;
    END
  END print_output[24]
  PIN print_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 796.000 361.010 800.000 ;
    END
  END print_output[25]
  PIN print_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END print_output[26]
  PIN print_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 346.840 800.000 347.440 ;
    END
  END print_output[27]
  PIN print_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END print_output[28]
  PIN print_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 53.080 800.000 53.680 ;
    END
  END print_output[29]
  PIN print_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END print_output[2]
  PIN print_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END print_output[30]
  PIN print_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END print_output[31]
  PIN print_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END print_output[3]
  PIN print_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 199.960 800.000 200.560 ;
    END
  END print_output[4]
  PIN print_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 796.000 708.770 800.000 ;
    END
  END print_output[5]
  PIN print_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 640.600 800.000 641.200 ;
    END
  END print_output[6]
  PIN print_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END print_output[7]
  PIN print_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END print_output[8]
  PIN print_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 334.600 800.000 335.200 ;
    END
  END print_output[9]
  PIN privilege_mode
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END privilege_mode
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 677.320 800.000 677.920 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 796.000 675.650 800.000 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 0.000 729.010 4.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 796.000 650.810 800.000 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 796.000 79.490 800.000 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 796.000 344.450 800.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 796.000 501.770 800.000 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 796.000 352.730 800.000 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 796.000 609.410 800.000 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 77.560 800.000 78.160 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 554.920 800.000 555.520 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 530.440 800.000 531.040 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 796.000 576.290 800.000 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 796.000 568.010 800.000 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 796.000 87.770 800.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 796.000 203.690 800.000 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END read_interactive_value[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 796.000 13.250 800.000 ;
    END
  END reset
  PIN reset_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 297.880 800.000 298.480 ;
    END
  END reset_mem_req
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 796.115 790.755 ;
      LAYER met1 ;
        RECT 0.070 6.500 799.870 791.140 ;
      LAYER met2 ;
        RECT 0.100 795.720 4.410 796.690 ;
        RECT 5.250 795.720 12.690 796.690 ;
        RECT 13.530 795.720 20.970 796.690 ;
        RECT 21.810 795.720 29.250 796.690 ;
        RECT 30.090 795.720 37.530 796.690 ;
        RECT 38.370 795.720 45.810 796.690 ;
        RECT 46.650 795.720 54.090 796.690 ;
        RECT 54.930 795.720 62.370 796.690 ;
        RECT 63.210 795.720 70.650 796.690 ;
        RECT 71.490 795.720 78.930 796.690 ;
        RECT 79.770 795.720 87.210 796.690 ;
        RECT 88.050 795.720 95.490 796.690 ;
        RECT 96.330 795.720 103.770 796.690 ;
        RECT 104.610 795.720 112.050 796.690 ;
        RECT 112.890 795.720 120.330 796.690 ;
        RECT 121.170 795.720 128.610 796.690 ;
        RECT 129.450 795.720 136.890 796.690 ;
        RECT 137.730 795.720 145.170 796.690 ;
        RECT 146.010 795.720 153.450 796.690 ;
        RECT 154.290 795.720 161.730 796.690 ;
        RECT 162.570 795.720 170.010 796.690 ;
        RECT 170.850 795.720 178.290 796.690 ;
        RECT 179.130 795.720 186.570 796.690 ;
        RECT 187.410 795.720 194.850 796.690 ;
        RECT 195.690 795.720 203.130 796.690 ;
        RECT 203.970 795.720 211.410 796.690 ;
        RECT 212.250 795.720 219.690 796.690 ;
        RECT 220.530 795.720 227.970 796.690 ;
        RECT 228.810 795.720 236.250 796.690 ;
        RECT 237.090 795.720 244.530 796.690 ;
        RECT 245.370 795.720 252.810 796.690 ;
        RECT 253.650 795.720 261.090 796.690 ;
        RECT 261.930 795.720 269.370 796.690 ;
        RECT 270.210 795.720 277.650 796.690 ;
        RECT 278.490 795.720 285.930 796.690 ;
        RECT 286.770 795.720 294.210 796.690 ;
        RECT 295.050 795.720 302.490 796.690 ;
        RECT 303.330 795.720 310.770 796.690 ;
        RECT 311.610 795.720 319.050 796.690 ;
        RECT 319.890 795.720 327.330 796.690 ;
        RECT 328.170 795.720 335.610 796.690 ;
        RECT 336.450 795.720 343.890 796.690 ;
        RECT 344.730 795.720 352.170 796.690 ;
        RECT 353.010 795.720 360.450 796.690 ;
        RECT 361.290 795.720 368.730 796.690 ;
        RECT 369.570 795.720 377.010 796.690 ;
        RECT 377.850 795.720 385.290 796.690 ;
        RECT 386.130 795.720 393.570 796.690 ;
        RECT 394.410 795.720 401.850 796.690 ;
        RECT 402.690 795.720 410.130 796.690 ;
        RECT 410.970 795.720 418.410 796.690 ;
        RECT 419.250 795.720 426.690 796.690 ;
        RECT 427.530 795.720 434.970 796.690 ;
        RECT 435.810 795.720 443.250 796.690 ;
        RECT 444.090 795.720 451.530 796.690 ;
        RECT 452.370 795.720 459.810 796.690 ;
        RECT 460.650 795.720 468.090 796.690 ;
        RECT 468.930 795.720 476.370 796.690 ;
        RECT 477.210 795.720 484.650 796.690 ;
        RECT 485.490 795.720 492.930 796.690 ;
        RECT 493.770 795.720 501.210 796.690 ;
        RECT 502.050 795.720 509.490 796.690 ;
        RECT 510.330 795.720 517.770 796.690 ;
        RECT 518.610 795.720 526.050 796.690 ;
        RECT 526.890 795.720 534.330 796.690 ;
        RECT 535.170 795.720 542.610 796.690 ;
        RECT 543.450 795.720 550.890 796.690 ;
        RECT 551.730 795.720 559.170 796.690 ;
        RECT 560.010 795.720 567.450 796.690 ;
        RECT 568.290 795.720 575.730 796.690 ;
        RECT 576.570 795.720 584.010 796.690 ;
        RECT 584.850 795.720 592.290 796.690 ;
        RECT 593.130 795.720 600.570 796.690 ;
        RECT 601.410 795.720 608.850 796.690 ;
        RECT 609.690 795.720 617.130 796.690 ;
        RECT 617.970 795.720 625.410 796.690 ;
        RECT 626.250 795.720 633.690 796.690 ;
        RECT 634.530 795.720 641.970 796.690 ;
        RECT 642.810 795.720 650.250 796.690 ;
        RECT 651.090 795.720 658.530 796.690 ;
        RECT 659.370 795.720 666.810 796.690 ;
        RECT 667.650 795.720 675.090 796.690 ;
        RECT 675.930 795.720 683.370 796.690 ;
        RECT 684.210 795.720 691.650 796.690 ;
        RECT 692.490 795.720 699.930 796.690 ;
        RECT 700.770 795.720 708.210 796.690 ;
        RECT 709.050 795.720 716.490 796.690 ;
        RECT 717.330 795.720 724.770 796.690 ;
        RECT 725.610 795.720 733.050 796.690 ;
        RECT 733.890 795.720 741.330 796.690 ;
        RECT 742.170 795.720 749.610 796.690 ;
        RECT 750.450 795.720 757.890 796.690 ;
        RECT 758.730 795.720 766.170 796.690 ;
        RECT 767.010 795.720 774.450 796.690 ;
        RECT 775.290 795.720 782.730 796.690 ;
        RECT 783.570 795.720 791.010 796.690 ;
        RECT 791.850 795.720 799.290 796.690 ;
        RECT 0.100 4.280 799.840 795.720 ;
        RECT 0.650 3.670 8.090 4.280 ;
        RECT 8.930 3.670 16.370 4.280 ;
        RECT 17.210 3.670 24.650 4.280 ;
        RECT 25.490 3.670 32.930 4.280 ;
        RECT 33.770 3.670 41.210 4.280 ;
        RECT 42.050 3.670 49.490 4.280 ;
        RECT 50.330 3.670 57.770 4.280 ;
        RECT 58.610 3.670 66.050 4.280 ;
        RECT 66.890 3.670 74.330 4.280 ;
        RECT 75.170 3.670 82.610 4.280 ;
        RECT 83.450 3.670 90.890 4.280 ;
        RECT 91.730 3.670 99.170 4.280 ;
        RECT 100.010 3.670 107.450 4.280 ;
        RECT 108.290 3.670 115.730 4.280 ;
        RECT 116.570 3.670 124.010 4.280 ;
        RECT 124.850 3.670 132.290 4.280 ;
        RECT 133.130 3.670 140.570 4.280 ;
        RECT 141.410 3.670 148.850 4.280 ;
        RECT 149.690 3.670 157.130 4.280 ;
        RECT 157.970 3.670 165.410 4.280 ;
        RECT 166.250 3.670 173.690 4.280 ;
        RECT 174.530 3.670 181.970 4.280 ;
        RECT 182.810 3.670 190.250 4.280 ;
        RECT 191.090 3.670 198.530 4.280 ;
        RECT 199.370 3.670 206.810 4.280 ;
        RECT 207.650 3.670 215.090 4.280 ;
        RECT 215.930 3.670 223.370 4.280 ;
        RECT 224.210 3.670 231.650 4.280 ;
        RECT 232.490 3.670 239.930 4.280 ;
        RECT 240.770 3.670 248.210 4.280 ;
        RECT 249.050 3.670 256.490 4.280 ;
        RECT 257.330 3.670 264.770 4.280 ;
        RECT 265.610 3.670 273.050 4.280 ;
        RECT 273.890 3.670 281.330 4.280 ;
        RECT 282.170 3.670 289.610 4.280 ;
        RECT 290.450 3.670 297.890 4.280 ;
        RECT 298.730 3.670 306.170 4.280 ;
        RECT 307.010 3.670 314.450 4.280 ;
        RECT 315.290 3.670 322.730 4.280 ;
        RECT 323.570 3.670 331.010 4.280 ;
        RECT 331.850 3.670 339.290 4.280 ;
        RECT 340.130 3.670 347.570 4.280 ;
        RECT 348.410 3.670 355.850 4.280 ;
        RECT 356.690 3.670 364.130 4.280 ;
        RECT 364.970 3.670 372.410 4.280 ;
        RECT 373.250 3.670 380.690 4.280 ;
        RECT 381.530 3.670 388.970 4.280 ;
        RECT 389.810 3.670 397.250 4.280 ;
        RECT 398.090 3.670 405.530 4.280 ;
        RECT 406.370 3.670 413.810 4.280 ;
        RECT 414.650 3.670 422.090 4.280 ;
        RECT 422.930 3.670 430.370 4.280 ;
        RECT 431.210 3.670 438.650 4.280 ;
        RECT 439.490 3.670 446.930 4.280 ;
        RECT 447.770 3.670 455.210 4.280 ;
        RECT 456.050 3.670 463.490 4.280 ;
        RECT 464.330 3.670 471.770 4.280 ;
        RECT 472.610 3.670 480.050 4.280 ;
        RECT 480.890 3.670 488.330 4.280 ;
        RECT 489.170 3.670 496.610 4.280 ;
        RECT 497.450 3.670 504.890 4.280 ;
        RECT 505.730 3.670 513.170 4.280 ;
        RECT 514.010 3.670 521.450 4.280 ;
        RECT 522.290 3.670 529.730 4.280 ;
        RECT 530.570 3.670 538.010 4.280 ;
        RECT 538.850 3.670 546.290 4.280 ;
        RECT 547.130 3.670 554.570 4.280 ;
        RECT 555.410 3.670 562.850 4.280 ;
        RECT 563.690 3.670 571.130 4.280 ;
        RECT 571.970 3.670 579.410 4.280 ;
        RECT 580.250 3.670 587.690 4.280 ;
        RECT 588.530 3.670 595.970 4.280 ;
        RECT 596.810 3.670 604.250 4.280 ;
        RECT 605.090 3.670 612.530 4.280 ;
        RECT 613.370 3.670 620.810 4.280 ;
        RECT 621.650 3.670 629.090 4.280 ;
        RECT 629.930 3.670 637.370 4.280 ;
        RECT 638.210 3.670 645.650 4.280 ;
        RECT 646.490 3.670 653.930 4.280 ;
        RECT 654.770 3.670 662.210 4.280 ;
        RECT 663.050 3.670 670.490 4.280 ;
        RECT 671.330 3.670 678.770 4.280 ;
        RECT 679.610 3.670 687.050 4.280 ;
        RECT 687.890 3.670 695.330 4.280 ;
        RECT 696.170 3.670 703.610 4.280 ;
        RECT 704.450 3.670 711.890 4.280 ;
        RECT 712.730 3.670 720.170 4.280 ;
        RECT 721.010 3.670 728.450 4.280 ;
        RECT 729.290 3.670 736.730 4.280 ;
        RECT 737.570 3.670 745.010 4.280 ;
        RECT 745.850 3.670 753.290 4.280 ;
        RECT 754.130 3.670 761.570 4.280 ;
        RECT 762.410 3.670 769.850 4.280 ;
        RECT 770.690 3.670 778.130 4.280 ;
        RECT 778.970 3.670 786.410 4.280 ;
        RECT 787.250 3.670 794.690 4.280 ;
        RECT 795.530 3.670 799.840 4.280 ;
      LAYER met3 ;
        RECT 4.400 793.880 796.000 794.745 ;
        RECT 4.000 788.480 796.000 793.880 ;
        RECT 4.000 787.080 795.600 788.480 ;
        RECT 4.000 783.040 796.000 787.080 ;
        RECT 4.400 781.640 796.000 783.040 ;
        RECT 4.000 776.240 796.000 781.640 ;
        RECT 4.000 774.840 795.600 776.240 ;
        RECT 4.000 770.800 796.000 774.840 ;
        RECT 4.400 769.400 796.000 770.800 ;
        RECT 4.000 764.000 796.000 769.400 ;
        RECT 4.000 762.600 795.600 764.000 ;
        RECT 4.000 758.560 796.000 762.600 ;
        RECT 4.400 757.160 796.000 758.560 ;
        RECT 4.000 751.760 796.000 757.160 ;
        RECT 4.000 750.360 795.600 751.760 ;
        RECT 4.000 746.320 796.000 750.360 ;
        RECT 4.400 744.920 796.000 746.320 ;
        RECT 4.000 739.520 796.000 744.920 ;
        RECT 4.000 738.120 795.600 739.520 ;
        RECT 4.000 734.080 796.000 738.120 ;
        RECT 4.400 732.680 796.000 734.080 ;
        RECT 4.000 727.280 796.000 732.680 ;
        RECT 4.000 725.880 795.600 727.280 ;
        RECT 4.000 721.840 796.000 725.880 ;
        RECT 4.400 720.440 796.000 721.840 ;
        RECT 4.000 715.040 796.000 720.440 ;
        RECT 4.000 713.640 795.600 715.040 ;
        RECT 4.000 709.600 796.000 713.640 ;
        RECT 4.400 708.200 796.000 709.600 ;
        RECT 4.000 702.800 796.000 708.200 ;
        RECT 4.000 701.400 795.600 702.800 ;
        RECT 4.000 697.360 796.000 701.400 ;
        RECT 4.400 695.960 796.000 697.360 ;
        RECT 4.000 690.560 796.000 695.960 ;
        RECT 4.000 689.160 795.600 690.560 ;
        RECT 4.000 685.120 796.000 689.160 ;
        RECT 4.400 683.720 796.000 685.120 ;
        RECT 4.000 678.320 796.000 683.720 ;
        RECT 4.000 676.920 795.600 678.320 ;
        RECT 4.000 672.880 796.000 676.920 ;
        RECT 4.400 671.480 796.000 672.880 ;
        RECT 4.000 666.080 796.000 671.480 ;
        RECT 4.000 664.680 795.600 666.080 ;
        RECT 4.000 660.640 796.000 664.680 ;
        RECT 4.400 659.240 796.000 660.640 ;
        RECT 4.000 653.840 796.000 659.240 ;
        RECT 4.000 652.440 795.600 653.840 ;
        RECT 4.000 648.400 796.000 652.440 ;
        RECT 4.400 647.000 796.000 648.400 ;
        RECT 4.000 641.600 796.000 647.000 ;
        RECT 4.000 640.200 795.600 641.600 ;
        RECT 4.000 636.160 796.000 640.200 ;
        RECT 4.400 634.760 796.000 636.160 ;
        RECT 4.000 629.360 796.000 634.760 ;
        RECT 4.000 627.960 795.600 629.360 ;
        RECT 4.000 623.920 796.000 627.960 ;
        RECT 4.400 622.520 796.000 623.920 ;
        RECT 4.000 617.120 796.000 622.520 ;
        RECT 4.000 615.720 795.600 617.120 ;
        RECT 4.000 611.680 796.000 615.720 ;
        RECT 4.400 610.280 796.000 611.680 ;
        RECT 4.000 604.880 796.000 610.280 ;
        RECT 4.000 603.480 795.600 604.880 ;
        RECT 4.000 599.440 796.000 603.480 ;
        RECT 4.400 598.040 796.000 599.440 ;
        RECT 4.000 592.640 796.000 598.040 ;
        RECT 4.000 591.240 795.600 592.640 ;
        RECT 4.000 587.200 796.000 591.240 ;
        RECT 4.400 585.800 796.000 587.200 ;
        RECT 4.000 580.400 796.000 585.800 ;
        RECT 4.000 579.000 795.600 580.400 ;
        RECT 4.000 574.960 796.000 579.000 ;
        RECT 4.400 573.560 796.000 574.960 ;
        RECT 4.000 568.160 796.000 573.560 ;
        RECT 4.000 566.760 795.600 568.160 ;
        RECT 4.000 562.720 796.000 566.760 ;
        RECT 4.400 561.320 796.000 562.720 ;
        RECT 4.000 555.920 796.000 561.320 ;
        RECT 4.000 554.520 795.600 555.920 ;
        RECT 4.000 550.480 796.000 554.520 ;
        RECT 4.400 549.080 796.000 550.480 ;
        RECT 4.000 543.680 796.000 549.080 ;
        RECT 4.000 542.280 795.600 543.680 ;
        RECT 4.000 538.240 796.000 542.280 ;
        RECT 4.400 536.840 796.000 538.240 ;
        RECT 4.000 531.440 796.000 536.840 ;
        RECT 4.000 530.040 795.600 531.440 ;
        RECT 4.000 526.000 796.000 530.040 ;
        RECT 4.400 524.600 796.000 526.000 ;
        RECT 4.000 519.200 796.000 524.600 ;
        RECT 4.000 517.800 795.600 519.200 ;
        RECT 4.000 513.760 796.000 517.800 ;
        RECT 4.400 512.360 796.000 513.760 ;
        RECT 4.000 506.960 796.000 512.360 ;
        RECT 4.000 505.560 795.600 506.960 ;
        RECT 4.000 501.520 796.000 505.560 ;
        RECT 4.400 500.120 796.000 501.520 ;
        RECT 4.000 494.720 796.000 500.120 ;
        RECT 4.000 493.320 795.600 494.720 ;
        RECT 4.000 489.280 796.000 493.320 ;
        RECT 4.400 487.880 796.000 489.280 ;
        RECT 4.000 482.480 796.000 487.880 ;
        RECT 4.000 481.080 795.600 482.480 ;
        RECT 4.000 477.040 796.000 481.080 ;
        RECT 4.400 475.640 796.000 477.040 ;
        RECT 4.000 470.240 796.000 475.640 ;
        RECT 4.000 468.840 795.600 470.240 ;
        RECT 4.000 464.800 796.000 468.840 ;
        RECT 4.400 463.400 796.000 464.800 ;
        RECT 4.000 458.000 796.000 463.400 ;
        RECT 4.000 456.600 795.600 458.000 ;
        RECT 4.000 452.560 796.000 456.600 ;
        RECT 4.400 451.160 796.000 452.560 ;
        RECT 4.000 445.760 796.000 451.160 ;
        RECT 4.000 444.360 795.600 445.760 ;
        RECT 4.000 440.320 796.000 444.360 ;
        RECT 4.400 438.920 796.000 440.320 ;
        RECT 4.000 433.520 796.000 438.920 ;
        RECT 4.000 432.120 795.600 433.520 ;
        RECT 4.000 428.080 796.000 432.120 ;
        RECT 4.400 426.680 796.000 428.080 ;
        RECT 4.000 421.280 796.000 426.680 ;
        RECT 4.000 419.880 795.600 421.280 ;
        RECT 4.000 415.840 796.000 419.880 ;
        RECT 4.400 414.440 796.000 415.840 ;
        RECT 4.000 409.040 796.000 414.440 ;
        RECT 4.000 407.640 795.600 409.040 ;
        RECT 4.000 403.600 796.000 407.640 ;
        RECT 4.400 402.200 796.000 403.600 ;
        RECT 4.000 396.800 796.000 402.200 ;
        RECT 4.000 395.400 795.600 396.800 ;
        RECT 4.000 391.360 796.000 395.400 ;
        RECT 4.400 389.960 796.000 391.360 ;
        RECT 4.000 384.560 796.000 389.960 ;
        RECT 4.000 383.160 795.600 384.560 ;
        RECT 4.000 379.120 796.000 383.160 ;
        RECT 4.400 377.720 796.000 379.120 ;
        RECT 4.000 372.320 796.000 377.720 ;
        RECT 4.000 370.920 795.600 372.320 ;
        RECT 4.000 366.880 796.000 370.920 ;
        RECT 4.400 365.480 796.000 366.880 ;
        RECT 4.000 360.080 796.000 365.480 ;
        RECT 4.000 358.680 795.600 360.080 ;
        RECT 4.000 354.640 796.000 358.680 ;
        RECT 4.400 353.240 796.000 354.640 ;
        RECT 4.000 347.840 796.000 353.240 ;
        RECT 4.000 346.440 795.600 347.840 ;
        RECT 4.000 342.400 796.000 346.440 ;
        RECT 4.400 341.000 796.000 342.400 ;
        RECT 4.000 335.600 796.000 341.000 ;
        RECT 4.000 334.200 795.600 335.600 ;
        RECT 4.000 330.160 796.000 334.200 ;
        RECT 4.400 328.760 796.000 330.160 ;
        RECT 4.000 323.360 796.000 328.760 ;
        RECT 4.000 321.960 795.600 323.360 ;
        RECT 4.000 317.920 796.000 321.960 ;
        RECT 4.400 316.520 796.000 317.920 ;
        RECT 4.000 311.120 796.000 316.520 ;
        RECT 4.000 309.720 795.600 311.120 ;
        RECT 4.000 305.680 796.000 309.720 ;
        RECT 4.400 304.280 796.000 305.680 ;
        RECT 4.000 298.880 796.000 304.280 ;
        RECT 4.000 297.480 795.600 298.880 ;
        RECT 4.000 293.440 796.000 297.480 ;
        RECT 4.400 292.040 796.000 293.440 ;
        RECT 4.000 286.640 796.000 292.040 ;
        RECT 4.000 285.240 795.600 286.640 ;
        RECT 4.000 281.200 796.000 285.240 ;
        RECT 4.400 279.800 796.000 281.200 ;
        RECT 4.000 274.400 796.000 279.800 ;
        RECT 4.000 273.000 795.600 274.400 ;
        RECT 4.000 268.960 796.000 273.000 ;
        RECT 4.400 267.560 796.000 268.960 ;
        RECT 4.000 262.160 796.000 267.560 ;
        RECT 4.000 260.760 795.600 262.160 ;
        RECT 4.000 256.720 796.000 260.760 ;
        RECT 4.400 255.320 796.000 256.720 ;
        RECT 4.000 249.920 796.000 255.320 ;
        RECT 4.000 248.520 795.600 249.920 ;
        RECT 4.000 244.480 796.000 248.520 ;
        RECT 4.400 243.080 796.000 244.480 ;
        RECT 4.000 237.680 796.000 243.080 ;
        RECT 4.000 236.280 795.600 237.680 ;
        RECT 4.000 232.240 796.000 236.280 ;
        RECT 4.400 230.840 796.000 232.240 ;
        RECT 4.000 225.440 796.000 230.840 ;
        RECT 4.000 224.040 795.600 225.440 ;
        RECT 4.000 220.000 796.000 224.040 ;
        RECT 4.400 218.600 796.000 220.000 ;
        RECT 4.000 213.200 796.000 218.600 ;
        RECT 4.000 211.800 795.600 213.200 ;
        RECT 4.000 207.760 796.000 211.800 ;
        RECT 4.400 206.360 796.000 207.760 ;
        RECT 4.000 200.960 796.000 206.360 ;
        RECT 4.000 199.560 795.600 200.960 ;
        RECT 4.000 195.520 796.000 199.560 ;
        RECT 4.400 194.120 796.000 195.520 ;
        RECT 4.000 188.720 796.000 194.120 ;
        RECT 4.000 187.320 795.600 188.720 ;
        RECT 4.000 183.280 796.000 187.320 ;
        RECT 4.400 181.880 796.000 183.280 ;
        RECT 4.000 176.480 796.000 181.880 ;
        RECT 4.000 175.080 795.600 176.480 ;
        RECT 4.000 171.040 796.000 175.080 ;
        RECT 4.400 169.640 796.000 171.040 ;
        RECT 4.000 164.240 796.000 169.640 ;
        RECT 4.000 162.840 795.600 164.240 ;
        RECT 4.000 158.800 796.000 162.840 ;
        RECT 4.400 157.400 796.000 158.800 ;
        RECT 4.000 152.000 796.000 157.400 ;
        RECT 4.000 150.600 795.600 152.000 ;
        RECT 4.000 146.560 796.000 150.600 ;
        RECT 4.400 145.160 796.000 146.560 ;
        RECT 4.000 139.760 796.000 145.160 ;
        RECT 4.000 138.360 795.600 139.760 ;
        RECT 4.000 134.320 796.000 138.360 ;
        RECT 4.400 132.920 796.000 134.320 ;
        RECT 4.000 127.520 796.000 132.920 ;
        RECT 4.000 126.120 795.600 127.520 ;
        RECT 4.000 122.080 796.000 126.120 ;
        RECT 4.400 120.680 796.000 122.080 ;
        RECT 4.000 115.280 796.000 120.680 ;
        RECT 4.000 113.880 795.600 115.280 ;
        RECT 4.000 109.840 796.000 113.880 ;
        RECT 4.400 108.440 796.000 109.840 ;
        RECT 4.000 103.040 796.000 108.440 ;
        RECT 4.000 101.640 795.600 103.040 ;
        RECT 4.000 97.600 796.000 101.640 ;
        RECT 4.400 96.200 796.000 97.600 ;
        RECT 4.000 90.800 796.000 96.200 ;
        RECT 4.000 89.400 795.600 90.800 ;
        RECT 4.000 85.360 796.000 89.400 ;
        RECT 4.400 83.960 796.000 85.360 ;
        RECT 4.000 78.560 796.000 83.960 ;
        RECT 4.000 77.160 795.600 78.560 ;
        RECT 4.000 73.120 796.000 77.160 ;
        RECT 4.400 71.720 796.000 73.120 ;
        RECT 4.000 66.320 796.000 71.720 ;
        RECT 4.000 64.920 795.600 66.320 ;
        RECT 4.000 60.880 796.000 64.920 ;
        RECT 4.400 59.480 796.000 60.880 ;
        RECT 4.000 54.080 796.000 59.480 ;
        RECT 4.000 52.680 795.600 54.080 ;
        RECT 4.000 48.640 796.000 52.680 ;
        RECT 4.400 47.240 796.000 48.640 ;
        RECT 4.000 41.840 796.000 47.240 ;
        RECT 4.000 40.440 795.600 41.840 ;
        RECT 4.000 36.400 796.000 40.440 ;
        RECT 4.400 35.000 796.000 36.400 ;
        RECT 4.000 29.600 796.000 35.000 ;
        RECT 4.000 28.200 795.600 29.600 ;
        RECT 4.000 24.160 796.000 28.200 ;
        RECT 4.400 22.760 796.000 24.160 ;
        RECT 4.000 17.360 796.000 22.760 ;
        RECT 4.000 15.960 795.600 17.360 ;
        RECT 4.000 11.920 796.000 15.960 ;
        RECT 4.400 10.520 796.000 11.920 ;
        RECT 4.000 5.120 796.000 10.520 ;
        RECT 4.000 4.255 795.600 5.120 ;
      LAYER met4 ;
        RECT 46.295 11.735 97.440 787.265 ;
        RECT 99.840 11.735 174.240 787.265 ;
        RECT 176.640 11.735 251.040 787.265 ;
        RECT 253.440 11.735 327.840 787.265 ;
        RECT 330.240 11.735 404.640 787.265 ;
        RECT 407.040 11.735 481.440 787.265 ;
        RECT 483.840 11.735 558.240 787.265 ;
        RECT 560.640 11.735 635.040 787.265 ;
        RECT 637.440 11.735 695.225 787.265 ;
  END
END datapath
END LIBRARY

