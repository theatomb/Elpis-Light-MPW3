VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 1496.000 8.650 1500.000 ;
    END
  END clk
  PIN data_from_mem[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 7.520 1500.000 8.120 ;
    END
  END data_from_mem[0]
  PIN data_from_mem[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.650 1496.000 1281.930 1500.000 ;
    END
  END data_from_mem[100]
  PIN data_from_mem[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.670 1496.000 1298.950 1500.000 ;
    END
  END data_from_mem[101]
  PIN data_from_mem[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1207.040 1500.000 1207.640 ;
    END
  END data_from_mem[102]
  PIN data_from_mem[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1223.360 1500.000 1223.960 ;
    END
  END data_from_mem[103]
  PIN data_from_mem[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.010 0.000 1312.290 4.000 ;
    END
  END data_from_mem[104]
  PIN data_from_mem[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 1496.000 1316.430 1500.000 ;
    END
  END data_from_mem[105]
  PIN data_from_mem[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1334.200 4.000 1334.800 ;
    END
  END data_from_mem[106]
  PIN data_from_mem[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1254.640 1500.000 1255.240 ;
    END
  END data_from_mem[107]
  PIN data_from_mem[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1270.280 1500.000 1270.880 ;
    END
  END data_from_mem[108]
  PIN data_from_mem[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 1496.000 1368.870 1500.000 ;
    END
  END data_from_mem[109]
  PIN data_from_mem[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 1496.000 304.890 1500.000 ;
    END
  END data_from_mem[10]
  PIN data_from_mem[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.430 0.000 1393.710 4.000 ;
    END
  END data_from_mem[110]
  PIN data_from_mem[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1285.920 1500.000 1286.520 ;
    END
  END data_from_mem[111]
  PIN data_from_mem[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1317.880 1500.000 1318.480 ;
    END
  END data_from_mem[112]
  PIN data_from_mem[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END data_from_mem[113]
  PIN data_from_mem[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1349.160 1500.000 1349.760 ;
    END
  END data_from_mem[114]
  PIN data_from_mem[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1372.960 4.000 1373.560 ;
    END
  END data_from_mem[115]
  PIN data_from_mem[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.990 0.000 1410.270 4.000 ;
    END
  END data_from_mem[116]
  PIN data_from_mem[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1381.120 1500.000 1381.720 ;
    END
  END data_from_mem[117]
  PIN data_from_mem[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.720 4.000 1412.320 ;
    END
  END data_from_mem[118]
  PIN data_from_mem[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 0.000 1442.930 4.000 ;
    END
  END data_from_mem[119]
  PIN data_from_mem[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END data_from_mem[11]
  PIN data_from_mem[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.510 1496.000 1438.790 1500.000 ;
    END
  END data_from_mem[120]
  PIN data_from_mem[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 0.000 1459.030 4.000 ;
    END
  END data_from_mem[121]
  PIN data_from_mem[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 0.000 1475.590 4.000 ;
    END
  END data_from_mem[122]
  PIN data_from_mem[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.470 1496.000 1473.750 1500.000 ;
    END
  END data_from_mem[123]
  PIN data_from_mem[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1444.360 1500.000 1444.960 ;
    END
  END data_from_mem[124]
  PIN data_from_mem[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1460.000 1500.000 1460.600 ;
    END
  END data_from_mem[125]
  PIN data_from_mem[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 0.000 1491.690 4.000 ;
    END
  END data_from_mem[126]
  PIN data_from_mem[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1491.280 1500.000 1491.880 ;
    END
  END data_from_mem[127]
  PIN data_from_mem[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END data_from_mem[12]
  PIN data_from_mem[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 1496.000 409.770 1500.000 ;
    END
  END data_from_mem[13]
  PIN data_from_mem[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END data_from_mem[14]
  PIN data_from_mem[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 291.080 1500.000 291.680 ;
    END
  END data_from_mem[15]
  PIN data_from_mem[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 323.040 1500.000 323.640 ;
    END
  END data_from_mem[16]
  PIN data_from_mem[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END data_from_mem[17]
  PIN data_from_mem[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 1496.000 461.750 1500.000 ;
    END
  END data_from_mem[18]
  PIN data_from_mem[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 1496.000 496.710 1500.000 ;
    END
  END data_from_mem[19]
  PIN data_from_mem[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END data_from_mem[1]
  PIN data_from_mem[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 1496.000 514.190 1500.000 ;
    END
  END data_from_mem[20]
  PIN data_from_mem[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END data_from_mem[21]
  PIN data_from_mem[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 433.200 1500.000 433.800 ;
    END
  END data_from_mem[22]
  PIN data_from_mem[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END data_from_mem[23]
  PIN data_from_mem[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 1496.000 566.630 1500.000 ;
    END
  END data_from_mem[24]
  PIN data_from_mem[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 465.160 1500.000 465.760 ;
    END
  END data_from_mem[25]
  PIN data_from_mem[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 480.800 1500.000 481.400 ;
    END
  END data_from_mem[26]
  PIN data_from_mem[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 1496.000 619.070 1500.000 ;
    END
  END data_from_mem[27]
  PIN data_from_mem[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 1496.000 636.550 1500.000 ;
    END
  END data_from_mem[28]
  PIN data_from_mem[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 512.760 1500.000 513.360 ;
    END
  END data_from_mem[29]
  PIN data_from_mem[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END data_from_mem[2]
  PIN data_from_mem[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 528.400 1500.000 529.000 ;
    END
  END data_from_mem[30]
  PIN data_from_mem[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 559.680 1500.000 560.280 ;
    END
  END data_from_mem[31]
  PIN data_from_mem[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END data_from_mem[32]
  PIN data_from_mem[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END data_from_mem[33]
  PIN data_from_mem[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 607.280 1500.000 607.880 ;
    END
  END data_from_mem[34]
  PIN data_from_mem[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 622.920 1500.000 623.520 ;
    END
  END data_from_mem[35]
  PIN data_from_mem[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.120 4.000 769.720 ;
    END
  END data_from_mem[36]
  PIN data_from_mem[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 654.880 1500.000 655.480 ;
    END
  END data_from_mem[37]
  PIN data_from_mem[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 670.520 1500.000 671.120 ;
    END
  END data_from_mem[38]
  PIN data_from_mem[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.160 4.000 788.760 ;
    END
  END data_from_mem[39]
  PIN data_from_mem[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END data_from_mem[3]
  PIN data_from_mem[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 686.160 1500.000 686.760 ;
    END
  END data_from_mem[40]
  PIN data_from_mem[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 827.600 4.000 828.200 ;
    END
  END data_from_mem[41]
  PIN data_from_mem[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 0.000 806.750 4.000 ;
    END
  END data_from_mem[42]
  PIN data_from_mem[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 0.000 823.310 4.000 ;
    END
  END data_from_mem[43]
  PIN data_from_mem[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 0.000 839.410 4.000 ;
    END
  END data_from_mem[44]
  PIN data_from_mem[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 1496.000 775.930 1500.000 ;
    END
  END data_from_mem[45]
  PIN data_from_mem[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 717.440 1500.000 718.040 ;
    END
  END data_from_mem[46]
  PIN data_from_mem[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END data_from_mem[47]
  PIN data_from_mem[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 1496.000 793.410 1500.000 ;
    END
  END data_from_mem[48]
  PIN data_from_mem[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.080 4.000 886.680 ;
    END
  END data_from_mem[49]
  PIN data_from_mem[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END data_from_mem[4]
  PIN data_from_mem[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END data_from_mem[50]
  PIN data_from_mem[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 780.680 1500.000 781.280 ;
    END
  END data_from_mem[51]
  PIN data_from_mem[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END data_from_mem[52]
  PIN data_from_mem[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 1496.000 845.850 1500.000 ;
    END
  END data_from_mem[53]
  PIN data_from_mem[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.450 0.000 904.730 4.000 ;
    END
  END data_from_mem[54]
  PIN data_from_mem[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 828.280 1500.000 828.880 ;
    END
  END data_from_mem[55]
  PIN data_from_mem[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END data_from_mem[56]
  PIN data_from_mem[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 1496.000 897.830 1500.000 ;
    END
  END data_from_mem[57]
  PIN data_from_mem[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 843.920 1500.000 844.520 ;
    END
  END data_from_mem[58]
  PIN data_from_mem[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 859.560 1500.000 860.160 ;
    END
  END data_from_mem[59]
  PIN data_from_mem[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END data_from_mem[5]
  PIN data_from_mem[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 0.000 970.050 4.000 ;
    END
  END data_from_mem[60]
  PIN data_from_mem[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END data_from_mem[61]
  PIN data_from_mem[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 944.560 4.000 945.160 ;
    END
  END data_from_mem[62]
  PIN data_from_mem[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 963.600 4.000 964.200 ;
    END
  END data_from_mem[63]
  PIN data_from_mem[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 4.000 ;
    END
  END data_from_mem[64]
  PIN data_from_mem[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.530 0.000 1018.810 4.000 ;
    END
  END data_from_mem[65]
  PIN data_from_mem[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.090 0.000 1035.370 4.000 ;
    END
  END data_from_mem[66]
  PIN data_from_mem[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 939.120 1500.000 939.720 ;
    END
  END data_from_mem[67]
  PIN data_from_mem[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 1496.000 967.750 1500.000 ;
    END
  END data_from_mem[68]
  PIN data_from_mem[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 954.760 1500.000 955.360 ;
    END
  END data_from_mem[69]
  PIN data_from_mem[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END data_from_mem[6]
  PIN data_from_mem[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 970.400 1500.000 971.000 ;
    END
  END data_from_mem[70]
  PIN data_from_mem[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 0.000 1051.470 4.000 ;
    END
  END data_from_mem[71]
  PIN data_from_mem[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 1496.000 1002.710 1500.000 ;
    END
  END data_from_mem[72]
  PIN data_from_mem[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 0.000 1067.570 4.000 ;
    END
  END data_from_mem[73]
  PIN data_from_mem[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 1496.000 1037.670 1500.000 ;
    END
  END data_from_mem[74]
  PIN data_from_mem[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.800 4.000 1042.400 ;
    END
  END data_from_mem[75]
  PIN data_from_mem[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1033.640 1500.000 1034.240 ;
    END
  END data_from_mem[76]
  PIN data_from_mem[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1049.280 1500.000 1049.880 ;
    END
  END data_from_mem[77]
  PIN data_from_mem[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 0.000 1100.230 4.000 ;
    END
  END data_from_mem[78]
  PIN data_from_mem[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1080.560 4.000 1081.160 ;
    END
  END data_from_mem[79]
  PIN data_from_mem[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 165.280 1500.000 165.880 ;
    END
  END data_from_mem[7]
  PIN data_from_mem[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1100.280 4.000 1100.880 ;
    END
  END data_from_mem[80]
  PIN data_from_mem[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.040 4.000 1139.640 ;
    END
  END data_from_mem[81]
  PIN data_from_mem[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 0.000 1116.790 4.000 ;
    END
  END data_from_mem[82]
  PIN data_from_mem[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.350 1496.000 1072.630 1500.000 ;
    END
  END data_from_mem[83]
  PIN data_from_mem[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.270 0.000 1165.550 4.000 ;
    END
  END data_from_mem[84]
  PIN data_from_mem[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END data_from_mem[85]
  PIN data_from_mem[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.800 4.000 1178.400 ;
    END
  END data_from_mem[86]
  PIN data_from_mem[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1112.520 1500.000 1113.120 ;
    END
  END data_from_mem[87]
  PIN data_from_mem[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.240 4.000 1217.840 ;
    END
  END data_from_mem[88]
  PIN data_from_mem[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 1496.000 1107.130 1500.000 ;
    END
  END data_from_mem[89]
  PIN data_from_mem[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END data_from_mem[8]
  PIN data_from_mem[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.280 4.000 1236.880 ;
    END
  END data_from_mem[90]
  PIN data_from_mem[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.810 1496.000 1142.090 1500.000 ;
    END
  END data_from_mem[91]
  PIN data_from_mem[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.770 1496.000 1177.050 1500.000 ;
    END
  END data_from_mem[92]
  PIN data_from_mem[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1143.800 1500.000 1144.400 ;
    END
  END data_from_mem[93]
  PIN data_from_mem[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.730 1496.000 1212.010 1500.000 ;
    END
  END data_from_mem[94]
  PIN data_from_mem[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1175.760 1500.000 1176.360 ;
    END
  END data_from_mem[95]
  PIN data_from_mem[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.210 1496.000 1229.490 1500.000 ;
    END
  END data_from_mem[96]
  PIN data_from_mem[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 1496.000 1246.970 1500.000 ;
    END
  END data_from_mem[97]
  PIN data_from_mem[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 1496.000 1264.450 1500.000 ;
    END
  END data_from_mem[98]
  PIN data_from_mem[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.720 4.000 1276.320 ;
    END
  END data_from_mem[99]
  PIN data_from_mem[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 1496.000 287.410 1500.000 ;
    END
  END data_from_mem[9]
  PIN hex_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 1496.000 148.030 1500.000 ;
    END
  END hex_out[0]
  PIN hex_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 212.200 1500.000 212.800 ;
    END
  END hex_out[10]
  PIN hex_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 228.520 1500.000 229.120 ;
    END
  END hex_out[11]
  PIN hex_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 1496.000 357.330 1500.000 ;
    END
  END hex_out[12]
  PIN hex_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 1496.000 427.250 1500.000 ;
    END
  END hex_out[13]
  PIN hex_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END hex_out[14]
  PIN hex_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END hex_out[15]
  PIN hex_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 338.680 1500.000 339.280 ;
    END
  END hex_out[16]
  PIN hex_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END hex_out[17]
  PIN hex_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 401.920 1500.000 402.520 ;
    END
  END hex_out[18]
  PIN hex_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 417.560 1500.000 418.160 ;
    END
  END hex_out[19]
  PIN hex_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 23.160 1500.000 23.760 ;
    END
  END hex_out[1]
  PIN hex_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END hex_out[20]
  PIN hex_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END hex_out[21]
  PIN hex_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END hex_out[22]
  PIN hex_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END hex_out[23]
  PIN hex_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END hex_out[24]
  PIN hex_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END hex_out[25]
  PIN hex_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 1496.000 601.590 1500.000 ;
    END
  END hex_out[26]
  PIN hex_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 0.000 660.010 4.000 ;
    END
  END hex_out[27]
  PIN hex_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END hex_out[28]
  PIN hex_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END hex_out[29]
  PIN hex_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END hex_out[2]
  PIN hex_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END hex_out[30]
  PIN hex_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 0.000 741.890 4.000 ;
    END
  END hex_out[31]
  PIN hex_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 1496.000 200.470 1500.000 ;
    END
  END hex_out[3]
  PIN hex_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 54.440 1500.000 55.040 ;
    END
  END hex_out[4]
  PIN hex_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 86.400 1500.000 87.000 ;
    END
  END hex_out[5]
  PIN hex_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 133.320 1500.000 133.920 ;
    END
  END hex_out[6]
  PIN hex_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END hex_out[7]
  PIN hex_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END hex_out[8]
  PIN hex_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 196.560 1500.000 197.160 ;
    END
  END hex_out[9]
  PIN hex_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 1496.000 78.110 1500.000 ;
    END
  END hex_req
  PIN is_mem_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 1496.000 130.550 1500.000 ;
    END
  END is_mem_ready
  PIN is_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 1496.000 113.070 1500.000 ;
    END
  END is_mem_req
  PIN is_mem_req_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END is_mem_req_reset
  PIN is_memory_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END is_memory_we
  PIN is_print_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 1496.000 95.590 1500.000 ;
    END
  END is_print_done
  PIN mem_addr_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END mem_addr_out[0]
  PIN mem_addr_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END mem_addr_out[10]
  PIN mem_addr_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END mem_addr_out[11]
  PIN mem_addr_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 244.160 1500.000 244.760 ;
    END
  END mem_addr_out[12]
  PIN mem_addr_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END mem_addr_out[13]
  PIN mem_addr_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 275.440 1500.000 276.040 ;
    END
  END mem_addr_out[14]
  PIN mem_addr_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 307.400 1500.000 308.000 ;
    END
  END mem_addr_out[15]
  PIN mem_addr_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END mem_addr_out[16]
  PIN mem_addr_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 370.640 1500.000 371.240 ;
    END
  END mem_addr_out[17]
  PIN mem_addr_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 1496.000 479.230 1500.000 ;
    END
  END mem_addr_out[18]
  PIN mem_addr_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END mem_addr_out[19]
  PIN mem_addr_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 1496.000 182.990 1500.000 ;
    END
  END mem_addr_out[1]
  PIN mem_addr_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END mem_addr_out[2]
  PIN mem_addr_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 1496.000 217.950 1500.000 ;
    END
  END mem_addr_out[3]
  PIN mem_addr_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 70.080 1500.000 70.680 ;
    END
  END mem_addr_out[4]
  PIN mem_addr_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 102.040 1500.000 102.640 ;
    END
  END mem_addr_out[5]
  PIN mem_addr_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END mem_addr_out[6]
  PIN mem_addr_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 1496.000 269.930 1500.000 ;
    END
  END mem_addr_out[7]
  PIN mem_addr_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END mem_addr_out[8]
  PIN mem_addr_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END mem_addr_out[9]
  PIN mem_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 1496.000 165.510 1500.000 ;
    END
  END mem_data_out[0]
  PIN mem_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.910 0.000 1296.190 4.000 ;
    END
  END mem_data_out[100]
  PIN mem_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1294.760 4.000 1295.360 ;
    END
  END mem_data_out[101]
  PIN mem_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1314.480 4.000 1315.080 ;
    END
  END mem_data_out[102]
  PIN mem_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1239.000 1500.000 1239.600 ;
    END
  END mem_data_out[103]
  PIN mem_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.570 0.000 1328.850 4.000 ;
    END
  END mem_data_out[104]
  PIN mem_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 1496.000 1333.910 1500.000 ;
    END
  END mem_data_out[105]
  PIN mem_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.670 0.000 1344.950 4.000 ;
    END
  END mem_data_out[106]
  PIN mem_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 0.000 1361.050 4.000 ;
    END
  END mem_data_out[107]
  PIN mem_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.110 1496.000 1351.390 1500.000 ;
    END
  END mem_data_out[108]
  PIN mem_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.330 0.000 1377.610 4.000 ;
    END
  END mem_data_out[109]
  PIN mem_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END mem_data_out[10]
  PIN mem_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.070 1496.000 1386.350 1500.000 ;
    END
  END mem_data_out[110]
  PIN mem_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1302.240 1500.000 1302.840 ;
    END
  END mem_data_out[111]
  PIN mem_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.550 1496.000 1403.830 1500.000 ;
    END
  END mem_data_out[112]
  PIN mem_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1333.520 1500.000 1334.120 ;
    END
  END mem_data_out[113]
  PIN mem_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 1496.000 1421.310 1500.000 ;
    END
  END mem_data_out[114]
  PIN mem_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1365.480 1500.000 1366.080 ;
    END
  END mem_data_out[115]
  PIN mem_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.090 0.000 1426.370 4.000 ;
    END
  END mem_data_out[116]
  PIN mem_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.680 4.000 1393.280 ;
    END
  END mem_data_out[117]
  PIN mem_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1396.760 1500.000 1397.360 ;
    END
  END mem_data_out[118]
  PIN mem_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1412.400 1500.000 1413.000 ;
    END
  END mem_data_out[119]
  PIN mem_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 1496.000 322.370 1500.000 ;
    END
  END mem_data_out[11]
  PIN mem_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END mem_data_out[120]
  PIN mem_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1428.040 1500.000 1428.640 ;
    END
  END mem_data_out[121]
  PIN mem_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 1496.000 1456.270 1500.000 ;
    END
  END mem_data_out[122]
  PIN mem_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.160 4.000 1451.760 ;
    END
  END mem_data_out[123]
  PIN mem_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 1496.000 1491.230 1500.000 ;
    END
  END mem_data_out[124]
  PIN mem_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1470.200 4.000 1470.800 ;
    END
  END mem_data_out[125]
  PIN mem_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1475.640 1500.000 1476.240 ;
    END
  END mem_data_out[126]
  PIN mem_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.920 4.000 1490.520 ;
    END
  END mem_data_out[127]
  PIN mem_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 1496.000 374.810 1500.000 ;
    END
  END mem_data_out[12]
  PIN mem_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 259.800 1500.000 260.400 ;
    END
  END mem_data_out[13]
  PIN mem_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END mem_data_out[14]
  PIN mem_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END mem_data_out[15]
  PIN mem_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 354.320 1500.000 354.920 ;
    END
  END mem_data_out[16]
  PIN mem_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END mem_data_out[17]
  PIN mem_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 4.000 ;
    END
  END mem_data_out[18]
  PIN mem_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END mem_data_out[19]
  PIN mem_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END mem_data_out[1]
  PIN mem_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END mem_data_out[20]
  PIN mem_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 1496.000 531.670 1500.000 ;
    END
  END mem_data_out[21]
  PIN mem_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 1496.000 549.150 1500.000 ;
    END
  END mem_data_out[22]
  PIN mem_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END mem_data_out[23]
  PIN mem_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END mem_data_out[24]
  PIN mem_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 0.000 627.350 4.000 ;
    END
  END mem_data_out[25]
  PIN mem_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 4.000 594.280 ;
    END
  END mem_data_out[26]
  PIN mem_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END mem_data_out[27]
  PIN mem_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END mem_data_out[28]
  PIN mem_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 1496.000 653.570 1500.000 ;
    END
  END mem_data_out[29]
  PIN mem_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END mem_data_out[2]
  PIN mem_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 1496.000 688.530 1500.000 ;
    END
  END mem_data_out[30]
  PIN mem_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END mem_data_out[31]
  PIN mem_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 575.320 1500.000 575.920 ;
    END
  END mem_data_out[32]
  PIN mem_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 591.640 1500.000 592.240 ;
    END
  END mem_data_out[33]
  PIN mem_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 0.000 757.990 4.000 ;
    END
  END mem_data_out[34]
  PIN mem_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END mem_data_out[35]
  PIN mem_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 638.560 1500.000 639.160 ;
    END
  END mem_data_out[36]
  PIN mem_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 0.000 774.090 4.000 ;
    END
  END mem_data_out[37]
  PIN mem_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 1496.000 706.010 1500.000 ;
    END
  END mem_data_out[38]
  PIN mem_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END mem_data_out[39]
  PIN mem_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 1496.000 234.970 1500.000 ;
    END
  END mem_data_out[3]
  PIN mem_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.370 0.000 790.650 4.000 ;
    END
  END mem_data_out[40]
  PIN mem_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 1496.000 723.490 1500.000 ;
    END
  END mem_data_out[41]
  PIN mem_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 1496.000 740.970 1500.000 ;
    END
  END mem_data_out[42]
  PIN mem_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END mem_data_out[43]
  PIN mem_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 1496.000 758.450 1500.000 ;
    END
  END mem_data_out[44]
  PIN mem_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 701.800 1500.000 702.400 ;
    END
  END mem_data_out[45]
  PIN mem_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END mem_data_out[46]
  PIN mem_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 733.760 1500.000 734.360 ;
    END
  END mem_data_out[47]
  PIN mem_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 749.400 1500.000 750.000 ;
    END
  END mem_data_out[48]
  PIN mem_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 1496.000 810.890 1500.000 ;
    END
  END mem_data_out[49]
  PIN mem_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END mem_data_out[4]
  PIN mem_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 765.040 1500.000 765.640 ;
    END
  END mem_data_out[50]
  PIN mem_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 797.000 1500.000 797.600 ;
    END
  END mem_data_out[51]
  PIN mem_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 1496.000 828.370 1500.000 ;
    END
  END mem_data_out[52]
  PIN mem_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 812.640 1500.000 813.240 ;
    END
  END mem_data_out[53]
  PIN mem_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 1496.000 863.330 1500.000 ;
    END
  END mem_data_out[54]
  PIN mem_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 0.000 920.830 4.000 ;
    END
  END mem_data_out[55]
  PIN mem_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.070 1496.000 880.350 1500.000 ;
    END
  END mem_data_out[56]
  PIN mem_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.120 4.000 905.720 ;
    END
  END mem_data_out[57]
  PIN mem_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END mem_data_out[58]
  PIN mem_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 875.880 1500.000 876.480 ;
    END
  END mem_data_out[59]
  PIN mem_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END mem_data_out[5]
  PIN mem_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.870 0.000 986.150 4.000 ;
    END
  END mem_data_out[60]
  PIN mem_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 891.520 1500.000 892.120 ;
    END
  END mem_data_out[61]
  PIN mem_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 1496.000 915.310 1500.000 ;
    END
  END mem_data_out[62]
  PIN mem_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 907.160 1500.000 907.760 ;
    END
  END mem_data_out[63]
  PIN mem_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 1496.000 932.790 1500.000 ;
    END
  END mem_data_out[64]
  PIN mem_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END mem_data_out[65]
  PIN mem_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 922.800 1500.000 923.400 ;
    END
  END mem_data_out[66]
  PIN mem_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 1496.000 950.270 1500.000 ;
    END
  END mem_data_out[67]
  PIN mem_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 1496.000 985.230 1500.000 ;
    END
  END mem_data_out[68]
  PIN mem_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END mem_data_out[69]
  PIN mem_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 148.960 1500.000 149.560 ;
    END
  END mem_data_out[6]
  PIN mem_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1022.080 4.000 1022.680 ;
    END
  END mem_data_out[70]
  PIN mem_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 986.040 1500.000 986.640 ;
    END
  END mem_data_out[71]
  PIN mem_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 1496.000 1020.190 1500.000 ;
    END
  END mem_data_out[72]
  PIN mem_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.850 0.000 1084.130 4.000 ;
    END
  END mem_data_out[73]
  PIN mem_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1001.680 1500.000 1002.280 ;
    END
  END mem_data_out[74]
  PIN mem_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1018.000 1500.000 1018.600 ;
    END
  END mem_data_out[75]
  PIN mem_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.870 1496.000 1055.150 1500.000 ;
    END
  END mem_data_out[76]
  PIN mem_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1064.920 1500.000 1065.520 ;
    END
  END mem_data_out[77]
  PIN mem_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1061.520 4.000 1062.120 ;
    END
  END mem_data_out[78]
  PIN mem_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1081.240 1500.000 1081.840 ;
    END
  END mem_data_out[79]
  PIN mem_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END mem_data_out[7]
  PIN mem_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.000 4.000 1120.600 ;
    END
  END mem_data_out[80]
  PIN mem_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1158.760 4.000 1159.360 ;
    END
  END mem_data_out[81]
  PIN mem_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.610 0.000 1132.890 4.000 ;
    END
  END mem_data_out[82]
  PIN mem_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.170 0.000 1149.450 4.000 ;
    END
  END mem_data_out[83]
  PIN mem_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 1496.000 1089.650 1500.000 ;
    END
  END mem_data_out[84]
  PIN mem_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1096.880 1500.000 1097.480 ;
    END
  END mem_data_out[85]
  PIN mem_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1197.520 4.000 1198.120 ;
    END
  END mem_data_out[86]
  PIN mem_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 0.000 1198.210 4.000 ;
    END
  END mem_data_out[87]
  PIN mem_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1128.160 1500.000 1128.760 ;
    END
  END mem_data_out[88]
  PIN mem_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.330 1496.000 1124.610 1500.000 ;
    END
  END mem_data_out[89]
  PIN mem_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END mem_data_out[8]
  PIN mem_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1256.000 4.000 1256.600 ;
    END
  END mem_data_out[90]
  PIN mem_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 1496.000 1159.570 1500.000 ;
    END
  END mem_data_out[91]
  PIN mem_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.250 1496.000 1194.530 1500.000 ;
    END
  END mem_data_out[92]
  PIN mem_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END mem_data_out[93]
  PIN mem_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1160.120 1500.000 1160.720 ;
    END
  END mem_data_out[94]
  PIN mem_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.590 0.000 1230.870 4.000 ;
    END
  END mem_data_out[95]
  PIN mem_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 0.000 1246.970 4.000 ;
    END
  END mem_data_out[96]
  PIN mem_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.250 0.000 1263.530 4.000 ;
    END
  END mem_data_out[97]
  PIN mem_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1191.400 1500.000 1192.000 ;
    END
  END mem_data_out[98]
  PIN mem_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.350 0.000 1279.630 4.000 ;
    END
  END mem_data_out[99]
  PIN mem_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END mem_data_out[9]
  PIN read_interactive_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 1496.000 43.150 1500.000 ;
    END
  END read_interactive_ready
  PIN read_interactive_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 1496.000 60.630 1500.000 ;
    END
  END read_interactive_req
  PIN read_interactive_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END read_interactive_value[0]
  PIN read_interactive_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END read_interactive_value[10]
  PIN read_interactive_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 1496.000 339.850 1500.000 ;
    END
  END read_interactive_value[11]
  PIN read_interactive_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 1496.000 392.290 1500.000 ;
    END
  END read_interactive_value[12]
  PIN read_interactive_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END read_interactive_value[13]
  PIN read_interactive_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END read_interactive_value[14]
  PIN read_interactive_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END read_interactive_value[15]
  PIN read_interactive_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 1496.000 444.270 1500.000 ;
    END
  END read_interactive_value[16]
  PIN read_interactive_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 386.280 1500.000 386.880 ;
    END
  END read_interactive_value[17]
  PIN read_interactive_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END read_interactive_value[18]
  PIN read_interactive_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 0.000 480.610 4.000 ;
    END
  END read_interactive_value[19]
  PIN read_interactive_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 38.800 1500.000 39.400 ;
    END
  END read_interactive_value[1]
  PIN read_interactive_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END read_interactive_value[20]
  PIN read_interactive_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END read_interactive_value[21]
  PIN read_interactive_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END read_interactive_value[22]
  PIN read_interactive_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 449.520 1500.000 450.120 ;
    END
  END read_interactive_value[23]
  PIN read_interactive_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 1496.000 584.110 1500.000 ;
    END
  END read_interactive_value[24]
  PIN read_interactive_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END read_interactive_value[25]
  PIN read_interactive_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 496.440 1500.000 497.040 ;
    END
  END read_interactive_value[26]
  PIN read_interactive_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END read_interactive_value[27]
  PIN read_interactive_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END read_interactive_value[28]
  PIN read_interactive_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 1496.000 671.050 1500.000 ;
    END
  END read_interactive_value[29]
  PIN read_interactive_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END read_interactive_value[2]
  PIN read_interactive_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 544.040 1500.000 544.640 ;
    END
  END read_interactive_value[30]
  PIN read_interactive_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END read_interactive_value[31]
  PIN read_interactive_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 1496.000 252.450 1500.000 ;
    END
  END read_interactive_value[3]
  PIN read_interactive_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END read_interactive_value[4]
  PIN read_interactive_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 117.680 1500.000 118.280 ;
    END
  END read_interactive_value[5]
  PIN read_interactive_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END read_interactive_value[6]
  PIN read_interactive_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END read_interactive_value[7]
  PIN read_interactive_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 180.920 1500.000 181.520 ;
    END
  END read_interactive_value[8]
  PIN read_interactive_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END read_interactive_value[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 1496.000 25.670 1500.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 1494.080 1488.480 ;
      LAYER met2 ;
        RECT 6.530 1495.720 8.090 1496.410 ;
        RECT 8.930 1495.720 25.110 1496.410 ;
        RECT 25.950 1495.720 42.590 1496.410 ;
        RECT 43.430 1495.720 60.070 1496.410 ;
        RECT 60.910 1495.720 77.550 1496.410 ;
        RECT 78.390 1495.720 95.030 1496.410 ;
        RECT 95.870 1495.720 112.510 1496.410 ;
        RECT 113.350 1495.720 129.990 1496.410 ;
        RECT 130.830 1495.720 147.470 1496.410 ;
        RECT 148.310 1495.720 164.950 1496.410 ;
        RECT 165.790 1495.720 182.430 1496.410 ;
        RECT 183.270 1495.720 199.910 1496.410 ;
        RECT 200.750 1495.720 217.390 1496.410 ;
        RECT 218.230 1495.720 234.410 1496.410 ;
        RECT 235.250 1495.720 251.890 1496.410 ;
        RECT 252.730 1495.720 269.370 1496.410 ;
        RECT 270.210 1495.720 286.850 1496.410 ;
        RECT 287.690 1495.720 304.330 1496.410 ;
        RECT 305.170 1495.720 321.810 1496.410 ;
        RECT 322.650 1495.720 339.290 1496.410 ;
        RECT 340.130 1495.720 356.770 1496.410 ;
        RECT 357.610 1495.720 374.250 1496.410 ;
        RECT 375.090 1495.720 391.730 1496.410 ;
        RECT 392.570 1495.720 409.210 1496.410 ;
        RECT 410.050 1495.720 426.690 1496.410 ;
        RECT 427.530 1495.720 443.710 1496.410 ;
        RECT 444.550 1495.720 461.190 1496.410 ;
        RECT 462.030 1495.720 478.670 1496.410 ;
        RECT 479.510 1495.720 496.150 1496.410 ;
        RECT 496.990 1495.720 513.630 1496.410 ;
        RECT 514.470 1495.720 531.110 1496.410 ;
        RECT 531.950 1495.720 548.590 1496.410 ;
        RECT 549.430 1495.720 566.070 1496.410 ;
        RECT 566.910 1495.720 583.550 1496.410 ;
        RECT 584.390 1495.720 601.030 1496.410 ;
        RECT 601.870 1495.720 618.510 1496.410 ;
        RECT 619.350 1495.720 635.990 1496.410 ;
        RECT 636.830 1495.720 653.010 1496.410 ;
        RECT 653.850 1495.720 670.490 1496.410 ;
        RECT 671.330 1495.720 687.970 1496.410 ;
        RECT 688.810 1495.720 705.450 1496.410 ;
        RECT 706.290 1495.720 722.930 1496.410 ;
        RECT 723.770 1495.720 740.410 1496.410 ;
        RECT 741.250 1495.720 757.890 1496.410 ;
        RECT 758.730 1495.720 775.370 1496.410 ;
        RECT 776.210 1495.720 792.850 1496.410 ;
        RECT 793.690 1495.720 810.330 1496.410 ;
        RECT 811.170 1495.720 827.810 1496.410 ;
        RECT 828.650 1495.720 845.290 1496.410 ;
        RECT 846.130 1495.720 862.770 1496.410 ;
        RECT 863.610 1495.720 879.790 1496.410 ;
        RECT 880.630 1495.720 897.270 1496.410 ;
        RECT 898.110 1495.720 914.750 1496.410 ;
        RECT 915.590 1495.720 932.230 1496.410 ;
        RECT 933.070 1495.720 949.710 1496.410 ;
        RECT 950.550 1495.720 967.190 1496.410 ;
        RECT 968.030 1495.720 984.670 1496.410 ;
        RECT 985.510 1495.720 1002.150 1496.410 ;
        RECT 1002.990 1495.720 1019.630 1496.410 ;
        RECT 1020.470 1495.720 1037.110 1496.410 ;
        RECT 1037.950 1495.720 1054.590 1496.410 ;
        RECT 1055.430 1495.720 1072.070 1496.410 ;
        RECT 1072.910 1495.720 1089.090 1496.410 ;
        RECT 1089.930 1495.720 1106.570 1496.410 ;
        RECT 1107.410 1495.720 1124.050 1496.410 ;
        RECT 1124.890 1495.720 1141.530 1496.410 ;
        RECT 1142.370 1495.720 1159.010 1496.410 ;
        RECT 1159.850 1495.720 1176.490 1496.410 ;
        RECT 1177.330 1495.720 1193.970 1496.410 ;
        RECT 1194.810 1495.720 1211.450 1496.410 ;
        RECT 1212.290 1495.720 1228.930 1496.410 ;
        RECT 1229.770 1495.720 1246.410 1496.410 ;
        RECT 1247.250 1495.720 1263.890 1496.410 ;
        RECT 1264.730 1495.720 1281.370 1496.410 ;
        RECT 1282.210 1495.720 1298.390 1496.410 ;
        RECT 1299.230 1495.720 1315.870 1496.410 ;
        RECT 1316.710 1495.720 1333.350 1496.410 ;
        RECT 1334.190 1495.720 1350.830 1496.410 ;
        RECT 1351.670 1495.720 1368.310 1496.410 ;
        RECT 1369.150 1495.720 1385.790 1496.410 ;
        RECT 1386.630 1495.720 1403.270 1496.410 ;
        RECT 1404.110 1495.720 1420.750 1496.410 ;
        RECT 1421.590 1495.720 1438.230 1496.410 ;
        RECT 1439.070 1495.720 1455.710 1496.410 ;
        RECT 1456.550 1495.720 1473.190 1496.410 ;
        RECT 1474.030 1495.720 1490.670 1496.410 ;
        RECT 1491.510 1495.720 1491.680 1496.410 ;
        RECT 6.530 4.280 1491.680 1495.720 ;
        RECT 6.530 3.670 7.630 4.280 ;
        RECT 8.470 3.670 23.730 4.280 ;
        RECT 24.570 3.670 39.830 4.280 ;
        RECT 40.670 3.670 56.390 4.280 ;
        RECT 57.230 3.670 72.490 4.280 ;
        RECT 73.330 3.670 89.050 4.280 ;
        RECT 89.890 3.670 105.150 4.280 ;
        RECT 105.990 3.670 121.710 4.280 ;
        RECT 122.550 3.670 137.810 4.280 ;
        RECT 138.650 3.670 154.370 4.280 ;
        RECT 155.210 3.670 170.470 4.280 ;
        RECT 171.310 3.670 186.570 4.280 ;
        RECT 187.410 3.670 203.130 4.280 ;
        RECT 203.970 3.670 219.230 4.280 ;
        RECT 220.070 3.670 235.790 4.280 ;
        RECT 236.630 3.670 251.890 4.280 ;
        RECT 252.730 3.670 268.450 4.280 ;
        RECT 269.290 3.670 284.550 4.280 ;
        RECT 285.390 3.670 301.110 4.280 ;
        RECT 301.950 3.670 317.210 4.280 ;
        RECT 318.050 3.670 333.310 4.280 ;
        RECT 334.150 3.670 349.870 4.280 ;
        RECT 350.710 3.670 365.970 4.280 ;
        RECT 366.810 3.670 382.530 4.280 ;
        RECT 383.370 3.670 398.630 4.280 ;
        RECT 399.470 3.670 415.190 4.280 ;
        RECT 416.030 3.670 431.290 4.280 ;
        RECT 432.130 3.670 447.850 4.280 ;
        RECT 448.690 3.670 463.950 4.280 ;
        RECT 464.790 3.670 480.050 4.280 ;
        RECT 480.890 3.670 496.610 4.280 ;
        RECT 497.450 3.670 512.710 4.280 ;
        RECT 513.550 3.670 529.270 4.280 ;
        RECT 530.110 3.670 545.370 4.280 ;
        RECT 546.210 3.670 561.930 4.280 ;
        RECT 562.770 3.670 578.030 4.280 ;
        RECT 578.870 3.670 594.590 4.280 ;
        RECT 595.430 3.670 610.690 4.280 ;
        RECT 611.530 3.670 626.790 4.280 ;
        RECT 627.630 3.670 643.350 4.280 ;
        RECT 644.190 3.670 659.450 4.280 ;
        RECT 660.290 3.670 676.010 4.280 ;
        RECT 676.850 3.670 692.110 4.280 ;
        RECT 692.950 3.670 708.670 4.280 ;
        RECT 709.510 3.670 724.770 4.280 ;
        RECT 725.610 3.670 741.330 4.280 ;
        RECT 742.170 3.670 757.430 4.280 ;
        RECT 758.270 3.670 773.530 4.280 ;
        RECT 774.370 3.670 790.090 4.280 ;
        RECT 790.930 3.670 806.190 4.280 ;
        RECT 807.030 3.670 822.750 4.280 ;
        RECT 823.590 3.670 838.850 4.280 ;
        RECT 839.690 3.670 855.410 4.280 ;
        RECT 856.250 3.670 871.510 4.280 ;
        RECT 872.350 3.670 888.070 4.280 ;
        RECT 888.910 3.670 904.170 4.280 ;
        RECT 905.010 3.670 920.270 4.280 ;
        RECT 921.110 3.670 936.830 4.280 ;
        RECT 937.670 3.670 952.930 4.280 ;
        RECT 953.770 3.670 969.490 4.280 ;
        RECT 970.330 3.670 985.590 4.280 ;
        RECT 986.430 3.670 1002.150 4.280 ;
        RECT 1002.990 3.670 1018.250 4.280 ;
        RECT 1019.090 3.670 1034.810 4.280 ;
        RECT 1035.650 3.670 1050.910 4.280 ;
        RECT 1051.750 3.670 1067.010 4.280 ;
        RECT 1067.850 3.670 1083.570 4.280 ;
        RECT 1084.410 3.670 1099.670 4.280 ;
        RECT 1100.510 3.670 1116.230 4.280 ;
        RECT 1117.070 3.670 1132.330 4.280 ;
        RECT 1133.170 3.670 1148.890 4.280 ;
        RECT 1149.730 3.670 1164.990 4.280 ;
        RECT 1165.830 3.670 1181.550 4.280 ;
        RECT 1182.390 3.670 1197.650 4.280 ;
        RECT 1198.490 3.670 1213.750 4.280 ;
        RECT 1214.590 3.670 1230.310 4.280 ;
        RECT 1231.150 3.670 1246.410 4.280 ;
        RECT 1247.250 3.670 1262.970 4.280 ;
        RECT 1263.810 3.670 1279.070 4.280 ;
        RECT 1279.910 3.670 1295.630 4.280 ;
        RECT 1296.470 3.670 1311.730 4.280 ;
        RECT 1312.570 3.670 1328.290 4.280 ;
        RECT 1329.130 3.670 1344.390 4.280 ;
        RECT 1345.230 3.670 1360.490 4.280 ;
        RECT 1361.330 3.670 1377.050 4.280 ;
        RECT 1377.890 3.670 1393.150 4.280 ;
        RECT 1393.990 3.670 1409.710 4.280 ;
        RECT 1410.550 3.670 1425.810 4.280 ;
        RECT 1426.650 3.670 1442.370 4.280 ;
        RECT 1443.210 3.670 1458.470 4.280 ;
        RECT 1459.310 3.670 1475.030 4.280 ;
        RECT 1475.870 3.670 1491.130 4.280 ;
      LAYER met3 ;
        RECT 4.000 1490.920 1495.600 1491.745 ;
        RECT 4.400 1490.880 1495.600 1490.920 ;
        RECT 4.400 1489.520 1496.000 1490.880 ;
        RECT 4.000 1476.640 1496.000 1489.520 ;
        RECT 4.000 1475.240 1495.600 1476.640 ;
        RECT 4.000 1471.200 1496.000 1475.240 ;
        RECT 4.400 1469.800 1496.000 1471.200 ;
        RECT 4.000 1461.000 1496.000 1469.800 ;
        RECT 4.000 1459.600 1495.600 1461.000 ;
        RECT 4.000 1452.160 1496.000 1459.600 ;
        RECT 4.400 1450.760 1496.000 1452.160 ;
        RECT 4.000 1445.360 1496.000 1450.760 ;
        RECT 4.000 1443.960 1495.600 1445.360 ;
        RECT 4.000 1432.440 1496.000 1443.960 ;
        RECT 4.400 1431.040 1496.000 1432.440 ;
        RECT 4.000 1429.040 1496.000 1431.040 ;
        RECT 4.000 1427.640 1495.600 1429.040 ;
        RECT 4.000 1413.400 1496.000 1427.640 ;
        RECT 4.000 1412.720 1495.600 1413.400 ;
        RECT 4.400 1412.000 1495.600 1412.720 ;
        RECT 4.400 1411.320 1496.000 1412.000 ;
        RECT 4.000 1397.760 1496.000 1411.320 ;
        RECT 4.000 1396.360 1495.600 1397.760 ;
        RECT 4.000 1393.680 1496.000 1396.360 ;
        RECT 4.400 1392.280 1496.000 1393.680 ;
        RECT 4.000 1382.120 1496.000 1392.280 ;
        RECT 4.000 1380.720 1495.600 1382.120 ;
        RECT 4.000 1373.960 1496.000 1380.720 ;
        RECT 4.400 1372.560 1496.000 1373.960 ;
        RECT 4.000 1366.480 1496.000 1372.560 ;
        RECT 4.000 1365.080 1495.600 1366.480 ;
        RECT 4.000 1354.240 1496.000 1365.080 ;
        RECT 4.400 1352.840 1496.000 1354.240 ;
        RECT 4.000 1350.160 1496.000 1352.840 ;
        RECT 4.000 1348.760 1495.600 1350.160 ;
        RECT 4.000 1335.200 1496.000 1348.760 ;
        RECT 4.400 1334.520 1496.000 1335.200 ;
        RECT 4.400 1333.800 1495.600 1334.520 ;
        RECT 4.000 1333.120 1495.600 1333.800 ;
        RECT 4.000 1318.880 1496.000 1333.120 ;
        RECT 4.000 1317.480 1495.600 1318.880 ;
        RECT 4.000 1315.480 1496.000 1317.480 ;
        RECT 4.400 1314.080 1496.000 1315.480 ;
        RECT 4.000 1303.240 1496.000 1314.080 ;
        RECT 4.000 1301.840 1495.600 1303.240 ;
        RECT 4.000 1295.760 1496.000 1301.840 ;
        RECT 4.400 1294.360 1496.000 1295.760 ;
        RECT 4.000 1286.920 1496.000 1294.360 ;
        RECT 4.000 1285.520 1495.600 1286.920 ;
        RECT 4.000 1276.720 1496.000 1285.520 ;
        RECT 4.400 1275.320 1496.000 1276.720 ;
        RECT 4.000 1271.280 1496.000 1275.320 ;
        RECT 4.000 1269.880 1495.600 1271.280 ;
        RECT 4.000 1257.000 1496.000 1269.880 ;
        RECT 4.400 1255.640 1496.000 1257.000 ;
        RECT 4.400 1255.600 1495.600 1255.640 ;
        RECT 4.000 1254.240 1495.600 1255.600 ;
        RECT 4.000 1240.000 1496.000 1254.240 ;
        RECT 4.000 1238.600 1495.600 1240.000 ;
        RECT 4.000 1237.280 1496.000 1238.600 ;
        RECT 4.400 1235.880 1496.000 1237.280 ;
        RECT 4.000 1224.360 1496.000 1235.880 ;
        RECT 4.000 1222.960 1495.600 1224.360 ;
        RECT 4.000 1218.240 1496.000 1222.960 ;
        RECT 4.400 1216.840 1496.000 1218.240 ;
        RECT 4.000 1208.040 1496.000 1216.840 ;
        RECT 4.000 1206.640 1495.600 1208.040 ;
        RECT 4.000 1198.520 1496.000 1206.640 ;
        RECT 4.400 1197.120 1496.000 1198.520 ;
        RECT 4.000 1192.400 1496.000 1197.120 ;
        RECT 4.000 1191.000 1495.600 1192.400 ;
        RECT 4.000 1178.800 1496.000 1191.000 ;
        RECT 4.400 1177.400 1496.000 1178.800 ;
        RECT 4.000 1176.760 1496.000 1177.400 ;
        RECT 4.000 1175.360 1495.600 1176.760 ;
        RECT 4.000 1161.120 1496.000 1175.360 ;
        RECT 4.000 1159.760 1495.600 1161.120 ;
        RECT 4.400 1159.720 1495.600 1159.760 ;
        RECT 4.400 1158.360 1496.000 1159.720 ;
        RECT 4.000 1144.800 1496.000 1158.360 ;
        RECT 4.000 1143.400 1495.600 1144.800 ;
        RECT 4.000 1140.040 1496.000 1143.400 ;
        RECT 4.400 1138.640 1496.000 1140.040 ;
        RECT 4.000 1129.160 1496.000 1138.640 ;
        RECT 4.000 1127.760 1495.600 1129.160 ;
        RECT 4.000 1121.000 1496.000 1127.760 ;
        RECT 4.400 1119.600 1496.000 1121.000 ;
        RECT 4.000 1113.520 1496.000 1119.600 ;
        RECT 4.000 1112.120 1495.600 1113.520 ;
        RECT 4.000 1101.280 1496.000 1112.120 ;
        RECT 4.400 1099.880 1496.000 1101.280 ;
        RECT 4.000 1097.880 1496.000 1099.880 ;
        RECT 4.000 1096.480 1495.600 1097.880 ;
        RECT 4.000 1082.240 1496.000 1096.480 ;
        RECT 4.000 1081.560 1495.600 1082.240 ;
        RECT 4.400 1080.840 1495.600 1081.560 ;
        RECT 4.400 1080.160 1496.000 1080.840 ;
        RECT 4.000 1065.920 1496.000 1080.160 ;
        RECT 4.000 1064.520 1495.600 1065.920 ;
        RECT 4.000 1062.520 1496.000 1064.520 ;
        RECT 4.400 1061.120 1496.000 1062.520 ;
        RECT 4.000 1050.280 1496.000 1061.120 ;
        RECT 4.000 1048.880 1495.600 1050.280 ;
        RECT 4.000 1042.800 1496.000 1048.880 ;
        RECT 4.400 1041.400 1496.000 1042.800 ;
        RECT 4.000 1034.640 1496.000 1041.400 ;
        RECT 4.000 1033.240 1495.600 1034.640 ;
        RECT 4.000 1023.080 1496.000 1033.240 ;
        RECT 4.400 1021.680 1496.000 1023.080 ;
        RECT 4.000 1019.000 1496.000 1021.680 ;
        RECT 4.000 1017.600 1495.600 1019.000 ;
        RECT 4.000 1004.040 1496.000 1017.600 ;
        RECT 4.400 1002.680 1496.000 1004.040 ;
        RECT 4.400 1002.640 1495.600 1002.680 ;
        RECT 4.000 1001.280 1495.600 1002.640 ;
        RECT 4.000 987.040 1496.000 1001.280 ;
        RECT 4.000 985.640 1495.600 987.040 ;
        RECT 4.000 984.320 1496.000 985.640 ;
        RECT 4.400 982.920 1496.000 984.320 ;
        RECT 4.000 971.400 1496.000 982.920 ;
        RECT 4.000 970.000 1495.600 971.400 ;
        RECT 4.000 964.600 1496.000 970.000 ;
        RECT 4.400 963.200 1496.000 964.600 ;
        RECT 4.000 955.760 1496.000 963.200 ;
        RECT 4.000 954.360 1495.600 955.760 ;
        RECT 4.000 945.560 1496.000 954.360 ;
        RECT 4.400 944.160 1496.000 945.560 ;
        RECT 4.000 940.120 1496.000 944.160 ;
        RECT 4.000 938.720 1495.600 940.120 ;
        RECT 4.000 925.840 1496.000 938.720 ;
        RECT 4.400 924.440 1496.000 925.840 ;
        RECT 4.000 923.800 1496.000 924.440 ;
        RECT 4.000 922.400 1495.600 923.800 ;
        RECT 4.000 908.160 1496.000 922.400 ;
        RECT 4.000 906.760 1495.600 908.160 ;
        RECT 4.000 906.120 1496.000 906.760 ;
        RECT 4.400 904.720 1496.000 906.120 ;
        RECT 4.000 892.520 1496.000 904.720 ;
        RECT 4.000 891.120 1495.600 892.520 ;
        RECT 4.000 887.080 1496.000 891.120 ;
        RECT 4.400 885.680 1496.000 887.080 ;
        RECT 4.000 876.880 1496.000 885.680 ;
        RECT 4.000 875.480 1495.600 876.880 ;
        RECT 4.000 867.360 1496.000 875.480 ;
        RECT 4.400 865.960 1496.000 867.360 ;
        RECT 4.000 860.560 1496.000 865.960 ;
        RECT 4.000 859.160 1495.600 860.560 ;
        RECT 4.000 847.640 1496.000 859.160 ;
        RECT 4.400 846.240 1496.000 847.640 ;
        RECT 4.000 844.920 1496.000 846.240 ;
        RECT 4.000 843.520 1495.600 844.920 ;
        RECT 4.000 829.280 1496.000 843.520 ;
        RECT 4.000 828.600 1495.600 829.280 ;
        RECT 4.400 827.880 1495.600 828.600 ;
        RECT 4.400 827.200 1496.000 827.880 ;
        RECT 4.000 813.640 1496.000 827.200 ;
        RECT 4.000 812.240 1495.600 813.640 ;
        RECT 4.000 808.880 1496.000 812.240 ;
        RECT 4.400 807.480 1496.000 808.880 ;
        RECT 4.000 798.000 1496.000 807.480 ;
        RECT 4.000 796.600 1495.600 798.000 ;
        RECT 4.000 789.160 1496.000 796.600 ;
        RECT 4.400 787.760 1496.000 789.160 ;
        RECT 4.000 781.680 1496.000 787.760 ;
        RECT 4.000 780.280 1495.600 781.680 ;
        RECT 4.000 770.120 1496.000 780.280 ;
        RECT 4.400 768.720 1496.000 770.120 ;
        RECT 4.000 766.040 1496.000 768.720 ;
        RECT 4.000 764.640 1495.600 766.040 ;
        RECT 4.000 750.400 1496.000 764.640 ;
        RECT 4.400 749.000 1495.600 750.400 ;
        RECT 4.000 734.760 1496.000 749.000 ;
        RECT 4.000 733.360 1495.600 734.760 ;
        RECT 4.000 731.360 1496.000 733.360 ;
        RECT 4.400 729.960 1496.000 731.360 ;
        RECT 4.000 718.440 1496.000 729.960 ;
        RECT 4.000 717.040 1495.600 718.440 ;
        RECT 4.000 711.640 1496.000 717.040 ;
        RECT 4.400 710.240 1496.000 711.640 ;
        RECT 4.000 702.800 1496.000 710.240 ;
        RECT 4.000 701.400 1495.600 702.800 ;
        RECT 4.000 691.920 1496.000 701.400 ;
        RECT 4.400 690.520 1496.000 691.920 ;
        RECT 4.000 687.160 1496.000 690.520 ;
        RECT 4.000 685.760 1495.600 687.160 ;
        RECT 4.000 672.880 1496.000 685.760 ;
        RECT 4.400 671.520 1496.000 672.880 ;
        RECT 4.400 671.480 1495.600 671.520 ;
        RECT 4.000 670.120 1495.600 671.480 ;
        RECT 4.000 655.880 1496.000 670.120 ;
        RECT 4.000 654.480 1495.600 655.880 ;
        RECT 4.000 653.160 1496.000 654.480 ;
        RECT 4.400 651.760 1496.000 653.160 ;
        RECT 4.000 639.560 1496.000 651.760 ;
        RECT 4.000 638.160 1495.600 639.560 ;
        RECT 4.000 633.440 1496.000 638.160 ;
        RECT 4.400 632.040 1496.000 633.440 ;
        RECT 4.000 623.920 1496.000 632.040 ;
        RECT 4.000 622.520 1495.600 623.920 ;
        RECT 4.000 614.400 1496.000 622.520 ;
        RECT 4.400 613.000 1496.000 614.400 ;
        RECT 4.000 608.280 1496.000 613.000 ;
        RECT 4.000 606.880 1495.600 608.280 ;
        RECT 4.000 594.680 1496.000 606.880 ;
        RECT 4.400 593.280 1496.000 594.680 ;
        RECT 4.000 592.640 1496.000 593.280 ;
        RECT 4.000 591.240 1495.600 592.640 ;
        RECT 4.000 576.320 1496.000 591.240 ;
        RECT 4.000 574.960 1495.600 576.320 ;
        RECT 4.400 574.920 1495.600 574.960 ;
        RECT 4.400 573.560 1496.000 574.920 ;
        RECT 4.000 560.680 1496.000 573.560 ;
        RECT 4.000 559.280 1495.600 560.680 ;
        RECT 4.000 555.920 1496.000 559.280 ;
        RECT 4.400 554.520 1496.000 555.920 ;
        RECT 4.000 545.040 1496.000 554.520 ;
        RECT 4.000 543.640 1495.600 545.040 ;
        RECT 4.000 536.200 1496.000 543.640 ;
        RECT 4.400 534.800 1496.000 536.200 ;
        RECT 4.000 529.400 1496.000 534.800 ;
        RECT 4.000 528.000 1495.600 529.400 ;
        RECT 4.000 516.480 1496.000 528.000 ;
        RECT 4.400 515.080 1496.000 516.480 ;
        RECT 4.000 513.760 1496.000 515.080 ;
        RECT 4.000 512.360 1495.600 513.760 ;
        RECT 4.000 497.440 1496.000 512.360 ;
        RECT 4.400 496.040 1495.600 497.440 ;
        RECT 4.000 481.800 1496.000 496.040 ;
        RECT 4.000 480.400 1495.600 481.800 ;
        RECT 4.000 477.720 1496.000 480.400 ;
        RECT 4.400 476.320 1496.000 477.720 ;
        RECT 4.000 466.160 1496.000 476.320 ;
        RECT 4.000 464.760 1495.600 466.160 ;
        RECT 4.000 458.000 1496.000 464.760 ;
        RECT 4.400 456.600 1496.000 458.000 ;
        RECT 4.000 450.520 1496.000 456.600 ;
        RECT 4.000 449.120 1495.600 450.520 ;
        RECT 4.000 438.960 1496.000 449.120 ;
        RECT 4.400 437.560 1496.000 438.960 ;
        RECT 4.000 434.200 1496.000 437.560 ;
        RECT 4.000 432.800 1495.600 434.200 ;
        RECT 4.000 419.240 1496.000 432.800 ;
        RECT 4.400 418.560 1496.000 419.240 ;
        RECT 4.400 417.840 1495.600 418.560 ;
        RECT 4.000 417.160 1495.600 417.840 ;
        RECT 4.000 402.920 1496.000 417.160 ;
        RECT 4.000 401.520 1495.600 402.920 ;
        RECT 4.000 399.520 1496.000 401.520 ;
        RECT 4.400 398.120 1496.000 399.520 ;
        RECT 4.000 387.280 1496.000 398.120 ;
        RECT 4.000 385.880 1495.600 387.280 ;
        RECT 4.000 380.480 1496.000 385.880 ;
        RECT 4.400 379.080 1496.000 380.480 ;
        RECT 4.000 371.640 1496.000 379.080 ;
        RECT 4.000 370.240 1495.600 371.640 ;
        RECT 4.000 360.760 1496.000 370.240 ;
        RECT 4.400 359.360 1496.000 360.760 ;
        RECT 4.000 355.320 1496.000 359.360 ;
        RECT 4.000 353.920 1495.600 355.320 ;
        RECT 4.000 341.720 1496.000 353.920 ;
        RECT 4.400 340.320 1496.000 341.720 ;
        RECT 4.000 339.680 1496.000 340.320 ;
        RECT 4.000 338.280 1495.600 339.680 ;
        RECT 4.000 324.040 1496.000 338.280 ;
        RECT 4.000 322.640 1495.600 324.040 ;
        RECT 4.000 322.000 1496.000 322.640 ;
        RECT 4.400 320.600 1496.000 322.000 ;
        RECT 4.000 308.400 1496.000 320.600 ;
        RECT 4.000 307.000 1495.600 308.400 ;
        RECT 4.000 302.280 1496.000 307.000 ;
        RECT 4.400 300.880 1496.000 302.280 ;
        RECT 4.000 292.080 1496.000 300.880 ;
        RECT 4.000 290.680 1495.600 292.080 ;
        RECT 4.000 283.240 1496.000 290.680 ;
        RECT 4.400 281.840 1496.000 283.240 ;
        RECT 4.000 276.440 1496.000 281.840 ;
        RECT 4.000 275.040 1495.600 276.440 ;
        RECT 4.000 263.520 1496.000 275.040 ;
        RECT 4.400 262.120 1496.000 263.520 ;
        RECT 4.000 260.800 1496.000 262.120 ;
        RECT 4.000 259.400 1495.600 260.800 ;
        RECT 4.000 245.160 1496.000 259.400 ;
        RECT 4.000 243.800 1495.600 245.160 ;
        RECT 4.400 243.760 1495.600 243.800 ;
        RECT 4.400 242.400 1496.000 243.760 ;
        RECT 4.000 229.520 1496.000 242.400 ;
        RECT 4.000 228.120 1495.600 229.520 ;
        RECT 4.000 224.760 1496.000 228.120 ;
        RECT 4.400 223.360 1496.000 224.760 ;
        RECT 4.000 213.200 1496.000 223.360 ;
        RECT 4.000 211.800 1495.600 213.200 ;
        RECT 4.000 205.040 1496.000 211.800 ;
        RECT 4.400 203.640 1496.000 205.040 ;
        RECT 4.000 197.560 1496.000 203.640 ;
        RECT 4.000 196.160 1495.600 197.560 ;
        RECT 4.000 185.320 1496.000 196.160 ;
        RECT 4.400 183.920 1496.000 185.320 ;
        RECT 4.000 181.920 1496.000 183.920 ;
        RECT 4.000 180.520 1495.600 181.920 ;
        RECT 4.000 166.280 1496.000 180.520 ;
        RECT 4.400 164.880 1495.600 166.280 ;
        RECT 4.000 149.960 1496.000 164.880 ;
        RECT 4.000 148.560 1495.600 149.960 ;
        RECT 4.000 146.560 1496.000 148.560 ;
        RECT 4.400 145.160 1496.000 146.560 ;
        RECT 4.000 134.320 1496.000 145.160 ;
        RECT 4.000 132.920 1495.600 134.320 ;
        RECT 4.000 126.840 1496.000 132.920 ;
        RECT 4.400 125.440 1496.000 126.840 ;
        RECT 4.000 118.680 1496.000 125.440 ;
        RECT 4.000 117.280 1495.600 118.680 ;
        RECT 4.000 107.800 1496.000 117.280 ;
        RECT 4.400 106.400 1496.000 107.800 ;
        RECT 4.000 103.040 1496.000 106.400 ;
        RECT 4.000 101.640 1495.600 103.040 ;
        RECT 4.000 88.080 1496.000 101.640 ;
        RECT 4.400 87.400 1496.000 88.080 ;
        RECT 4.400 86.680 1495.600 87.400 ;
        RECT 4.000 86.000 1495.600 86.680 ;
        RECT 4.000 71.080 1496.000 86.000 ;
        RECT 4.000 69.680 1495.600 71.080 ;
        RECT 4.000 68.360 1496.000 69.680 ;
        RECT 4.400 66.960 1496.000 68.360 ;
        RECT 4.000 55.440 1496.000 66.960 ;
        RECT 4.000 54.040 1495.600 55.440 ;
        RECT 4.000 49.320 1496.000 54.040 ;
        RECT 4.400 47.920 1496.000 49.320 ;
        RECT 4.000 39.800 1496.000 47.920 ;
        RECT 4.000 38.400 1495.600 39.800 ;
        RECT 4.000 29.600 1496.000 38.400 ;
        RECT 4.400 28.200 1496.000 29.600 ;
        RECT 4.000 24.160 1496.000 28.200 ;
        RECT 4.000 22.760 1495.600 24.160 ;
        RECT 4.000 10.560 1496.000 22.760 ;
        RECT 4.400 9.160 1496.000 10.560 ;
        RECT 4.000 8.520 1496.000 9.160 ;
        RECT 4.000 7.655 1495.600 8.520 ;
      LAYER met4 ;
        RECT 290.095 17.855 327.840 1486.305 ;
        RECT 330.240 17.855 404.640 1486.305 ;
        RECT 407.040 17.855 481.440 1486.305 ;
        RECT 483.840 17.855 558.240 1486.305 ;
        RECT 560.640 17.855 635.040 1486.305 ;
        RECT 637.440 17.855 711.840 1486.305 ;
        RECT 714.240 17.855 788.640 1486.305 ;
        RECT 791.040 17.855 865.440 1486.305 ;
        RECT 867.840 17.855 942.240 1486.305 ;
        RECT 944.640 17.855 1018.145 1486.305 ;
  END
END core
END LIBRARY

